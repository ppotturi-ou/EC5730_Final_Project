module lcd_timing_controller		(
						iCLK, 				// LCD display clock
						iRST_n, 			// systen reset
						//LCD SIDE
						oHD,				// LCD Horizontal sync 
						oVD,				// LCD Vertical sync 	
						oDEN,				// LCD Data Enable
						oLCD_R,				// LCD Red color data 
						oLCD_G,             // LCD Green color data  
						oLCD_B,             // LCD Blue color data  
						iDISPLAY_MODE
						);
//============================================================================
// PARAMETER declarations
//============================================================================
parameter H_LINE = 1056;
parameter V_LINE = 525;
parameter Hsync_Blank = 216;
parameter Hsync_Front_Porch = 40;
parameter Vertical_Back_Porch = 75;
parameter Vertical_Front_Porch = 50;
parameter hres_limit = 80;
parameter vres_limit = 40;
parameter tres_limit = 100;
parameter hres_limit1 = 8;
parameter vres_limit1 = 4;
parameter tres_limit1 = 10000;
parameter tres_limit12= 40000;
//===========================================================================
// PORT declarations
//===========================================================================
input			iCLK;   
input			iRST_n;
output	[7:0] oLCD_R;		
output   [7:0]	oLCD_G;
output   [7:0]	oLCD_B;
output			oHD;
output			oVD;
output			oDEN;
input	[1:0]	iDISPLAY_MODE;	
//=============================================================================
// REG/WIRE declarations
//=============================================================================
integer pic_cnt = 99;
integer pic_cnt1 = 9;
integer pic_cnt2 = 9999;
integer pic_cnt3 = 99;
integer res_cnt = 0;
integer vres_cnt = 0;
integer res_cnt1 = 0;
integer vres_cnt1 = 0;
reg		[10:0]  x_cnt;  
//reg		[10:0]  pic_cnt; 
//reg		[10:0]  res_cnt;  
reg		[9:0]	y_cnt; 
wire	[7:0]	mred;
wire	[7:0]	mgreen;
wire	[7:0]	mblue; 
wire			display_area;
reg				mhd;
reg				mvd;
reg				mden;
reg				oHD;
reg				oVD;
reg				oDEN;
reg		[7:0]	oLCD_R;
reg		[7:0]	oLCD_G;	
reg		[7:0]	oLCD_B;	
wire	[1:0]	msel;
wire	[1:0]	mselx;	
wire	[1:0]	msel1;
wire	[1:0]	mselx1;	
reg		[7:0]	red_1;
reg 	[7:0]	green_1;
reg 	[7:0]	blue_1;
reg		[7:0]	red_2;
reg 	[7:0]	green_2;
reg 	[7:0]	blue_2;
reg		[7:0]	red_3;
reg 	[7:0]	green_3;
reg 	[7:0]	blue_3;
reg		[7:0]	red_4;
reg 	[7:0]	green_4;
reg 	[7:0]	blue_4;
reg 	[7:0]	graycnt;
reg 	[7:0]	graycnt1;
reg	[7:0]	pattern_data;

reg	[7:0]	pattern_data_B [0:99] = '{8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF,8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'h00, 8'h00, 8'hFF, 8'hFF};
reg	[7:0]	pattern_data_G [0:99] = '{8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A,8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h13, 8'h13, 8'h5A, 8'h5A};
reg	[7:0]	pattern_data_R [0:99] = '{8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4, 8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4,8'h00, 8'h00, 8'h01, 8'h01, 8'hFF, 8'hFF, 8'hD4, 8'hD4, 8'hA4, 8'hA4};

reg	[7:0]	pattern_data_R1 [0:39999] = '{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hFA, 8'hF8, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF8, 8'hFA, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF1, 8'hE7, 8'hE0, 8'hDB, 8'hDB, 8'hDC, 8'hDD, 8'hDD, 8'hDC, 8'hDB, 8'hDB, 8'hE0, 8'hE8, 8'hF1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hDF, 8'hC9, 8'hB9, 8'hAD, 8'hAE, 8'hB0, 8'hB1, 8'hB1, 8'hB0, 8'hAE, 8'hAD, 8'hB9, 8'hCA, 8'hDF, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC8, 8'hA5, 8'h88, 8'h74, 8'h76, 8'h7A, 8'h7B, 8'h7B, 8'h7A, 8'h76, 8'h74, 8'h88, 8'hA6, 8'hC8, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFA, 8'hF7, 8'hE8, 8'hB3, 8'h86, 8'h62, 8'h49, 8'h4B, 8'h50, 8'h52, 8'h52, 8'h50, 8'h4B, 8'h49, 8'h62, 8'h87, 8'hB3, 8'hE8, 8'hF7, 8'hFA, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hE6, 8'hDB, 8'hCE, 8'h9B, 8'h70, 8'h4E, 8'h36, 8'h38, 8'h3D, 8'h3F, 8'h3F, 8'h3D, 8'h38, 8'h36, 8'h4E, 8'h72, 8'h9B, 8'hCE, 8'hDB, 8'hE6, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'hC7, 8'hAD, 8'hA7, 8'h84, 8'h65, 8'h4E, 8'h3C, 8'h3F, 8'h42, 8'h44, 8'h44, 8'h42, 8'h3F, 8'h3C, 8'h4E, 8'h67, 8'h84, 8'hA7, 8'hAD, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hA0, 8'h74, 8'h79, 8'h6B, 8'h5F, 8'h55, 8'h4F, 8'h50, 8'h53, 8'h53, 8'h53, 8'h53, 8'h50, 8'h4F, 8'h55, 8'h5F, 8'h6B, 8'h79, 8'h74, 8'hA1, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF7, 8'hCF, 8'h80, 8'h49, 8'h55, 8'h58, 8'h5A, 8'h5C, 8'h5D, 8'h5F, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5F, 8'h5D, 8'h5C, 8'h5A, 8'h58, 8'h55, 8'h49, 8'h81, 8'hD1, 8'hF7, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'hDB, 8'hB6, 8'h6B, 8'h36, 8'h44, 8'h50, 8'h59, 8'h61, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h61, 8'h59, 8'h50, 8'h44, 8'h36, 8'h6B, 8'hB8, 8'hDB, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hAE, 8'h97, 8'h62, 8'h3C, 8'h48, 8'h53, 8'h5C, 8'h63, 8'h68, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h68, 8'h63, 8'h5C, 8'h53, 8'h48, 8'h3C, 8'h62, 8'h98, 8'hAE, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h76, 8'h72, 8'h5E, 8'h4F, 8'h56, 8'h5C, 8'h60, 8'h64, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h64, 8'h60, 8'h5C, 8'h56, 8'h4F, 8'h5E, 8'h72, 8'h76, 8'hB7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF7, 8'h9D, 8'h4B, 8'h56, 8'h5B, 8'h5D, 8'h60, 8'h63, 8'h64, 8'h65, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h65, 8'h64, 8'h63, 8'h60, 8'h5D, 8'h5B, 8'h56, 8'h4B, 8'h9D, 8'hF7, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hDB, 8'h86, 8'h38, 8'h49, 8'h5B, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h5A, 8'h49, 8'h38, 8'h86, 8'hDB, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'hAD, 8'h75, 8'h3E, 8'h4D, 8'h5E, 8'h68, 8'h68, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h68, 8'h68, 8'h5D, 8'h4D, 8'h3E, 8'h75, 8'hAD, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h74, 8'h64, 8'h50, 8'h59, 8'h61, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h61, 8'h58, 8'h50, 8'h64, 8'h74, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF7, 8'h91, 8'h49, 8'h58, 8'h5E, 8'h62, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h62, 8'h5E, 8'h58, 8'h49, 8'h91, 8'hF7, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hDB, 8'h7A, 8'h36, 8'h54, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h54, 8'h36, 8'h7A, 8'hDB, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'hAD, 8'h6D, 8'h3C, 8'h57, 8'h68, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h68, 8'h57, 8'h3C, 8'h6D, 8'hAD, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'h74, 8'h61, 8'h4F, 8'h5E, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h5E, 8'h4F, 8'h61, 8'h74, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hB5, 8'h49, 8'h59, 8'h5D, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h5D, 8'h59, 8'h49, 8'hB6, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'h9D, 8'h36, 8'h56, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h56, 8'h36, 8'h9D, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB9, 8'h84, 8'h3C, 8'h59, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h59, 8'h3C, 8'h84, 8'hB9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h88, 8'h69, 8'h4F, 8'h5F, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h5F, 8'h4F, 8'h69, 8'h88, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF7, 8'h62, 8'h55, 8'h5D, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h5D, 8'h54, 8'h62, 8'hF7, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hDB, 8'h4E, 8'h4C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4B, 8'h4E, 8'hDB, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hAD, 8'h4D, 8'h51, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h50, 8'h4D, 8'hAD, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'h75, 8'h54, 8'h5A, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5A, 8'h54, 8'h75, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hD7, 8'h4A, 8'h5B, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h62, 8'h5B, 8'h4A, 8'hD7, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hBC, 8'h36, 8'h5F, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5F, 8'h36, 8'hBC, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h98, 8'h3D, 8'h62, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h62, 8'h3D, 8'h98, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC1, 8'h6D, 8'h4F, 8'h64, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h64, 8'h4F, 8'h6D, 8'hC1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hAA, 8'h4D, 8'h5D, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5D, 8'h4D, 8'hAA, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h91, 8'h3F, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h3F, 8'h91, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h7A, 8'h45, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h45, 8'h7A, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h63, 8'h55, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h55, 8'h63, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h95, 8'h51, 8'h61, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h61, 8'h51, 8'h95, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'h7D, 8'h4A, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h4A, 8'h7D, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD3, 8'h6C, 8'h4F, 8'h69, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h69, 8'h4F, 8'h6C, 8'hD3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5D, 8'h5A, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h5A, 8'h5D, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h9A, 8'h51, 8'h62, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h62, 8'h51, 8'h99, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h81, 8'h4E, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4E, 8'h81, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'h6E, 8'h53, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h53, 8'h6E, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCB, 8'h5C, 8'h5C, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5C, 8'h5C, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hB5, 8'h4E, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h4F, 8'hB5, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h9B, 8'h4A, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4B, 8'h9B, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'h7F, 8'h50, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h50, 8'h7F, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'h61, 8'h59, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h68, 8'h69, 8'h69, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h69, 8'h69, 8'h68, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5A, 8'h61, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h4A, 8'h62, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h67, 8'h67, 8'h67, 8'h66, 8'h65, 8'h65, 8'h65, 8'h65, 8'h66, 8'h67, 8'h67, 8'h67, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h62, 8'h4A, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'h41, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h63, 8'h61, 8'h60, 8'h60, 8'h5E, 8'h5D, 8'h5E, 8'h5E, 8'h5E, 8'h5E, 8'h5D, 8'h5E, 8'h60, 8'h60, 8'h61, 8'h63, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h41, 8'hCD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA6, 8'h47, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h63, 8'h5D, 8'h59, 8'h55, 8'h53, 8'h50, 8'h4F, 8'h51, 8'h53, 8'h53, 8'h51, 8'h4F, 8'h50, 8'h53, 8'h55, 8'h59, 8'h5D, 8'h63, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h47, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h77, 8'h55, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h68, 8'h5F, 8'h56, 8'h4E, 8'h47, 8'h42, 8'h3E, 8'h3C, 8'h40, 8'h45, 8'h45, 8'h40, 8'h3C, 8'h3E, 8'h42, 8'h47, 8'h4E, 8'h56, 8'h5F, 8'h68, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h55, 8'h77, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'h52, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h5D, 8'h52, 8'h4B, 8'h43, 8'h3D, 8'h37, 8'h36, 8'h3B, 8'h41, 8'h41, 8'h3B, 8'h36, 8'h37, 8'h3D, 8'h43, 8'h4B, 8'h52, 8'h5D, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h52, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h40, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h60, 8'h5D, 8'h5B, 8'h58, 8'h57, 8'h54, 8'h50, 8'h4A, 8'h49, 8'h4E, 8'h55, 8'h55, 8'h4E, 8'h49, 8'h4A, 8'h50, 8'h54, 8'h57, 8'h58, 8'h5B, 8'h5D, 8'h60, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h40, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC7, 8'h43, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h5E, 8'h55, 8'h4F, 8'h5B, 8'h67, 8'h72, 8'h7A, 8'h7A, 8'h76, 8'h74, 8'h79, 8'h7E, 8'h7E, 8'h79, 8'h74, 8'h76, 8'h7A, 8'h7A, 8'h72, 8'h67, 8'h5B, 8'h4F, 8'h55, 8'h5E, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h43, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA0, 8'h4E, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h68, 8'h65, 8'h56, 8'h48, 8'h3D, 8'h5B, 8'h7B, 8'h96, 8'hAB, 8'hB0, 8'hAD, 8'hAD, 8'hAF, 8'hB2, 8'hB2, 8'hAF, 8'hAD, 8'hAD, 8'hB0, 8'hAB, 8'h95, 8'h7B, 8'h5A, 8'h3D, 8'h48, 8'h56, 8'h65, 8'h68, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4E, 8'hA0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h7F, 8'h58, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h63, 8'h53, 8'h43, 8'h36, 8'h61, 8'h8E, 8'hB4, 8'hD3, 8'hDC, 8'hDB, 8'hDB, 8'hDC, 8'hDD, 8'hDD, 8'hDC, 8'hDB, 8'hDB, 8'hDC, 8'hD3, 8'hB4, 8'h8E, 8'h60, 8'h36, 8'h43, 8'h53, 8'h63, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h58, 8'h7F, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h68, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h65, 8'h60, 8'h5D, 8'h59, 8'h55, 8'h4A, 8'h76, 8'hA5, 8'hCD, 8'hED, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF8, 8'hF8, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hED, 8'hCC, 8'hA5, 8'h75, 8'h4A, 8'h55, 8'h59, 8'h5D, 8'h60, 8'h65, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h68, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'h5B, 8'h62, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h61, 8'h55, 8'h52, 8'h67, 8'h7A, 8'h75, 8'h98, 8'hBE, 8'hDD, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hDC, 8'hBE, 8'h97, 8'h75, 8'h7A, 8'h67, 8'h52, 8'h55, 8'h62, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h62, 8'h5B, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'h52, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h69, 8'h5E, 8'h47, 8'h45, 8'h7A, 8'hA9, 8'hAD, 8'hC2, 8'hD8, 8'hEB, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hEB, 8'hD8, 8'hC2, 8'hAD, 8'hA9, 8'h7A, 8'h44, 8'h48, 8'h5E, 8'h69, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h52, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'h4C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h5B, 8'h42, 8'h42, 8'h8D, 8'hD1, 8'hDB, 8'hE4, 8'hEE, 8'hF6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF6, 8'hEE, 8'hE4, 8'hDB, 8'hD1, 8'h8D, 8'h41, 8'h43, 8'h5C, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4C, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'h4C, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h65, 8'h60, 8'h5A, 8'h53, 8'h55, 8'hA4, 8'hEB, 8'hF7, 8'hF9, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hF9, 8'hF7, 8'hEB, 8'hA4, 8'h55, 8'h53, 8'h5B, 8'h60, 8'h65, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4C, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAC, 8'h51, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h62, 8'h52, 8'h5C, 8'h77, 8'h7E, 8'hBC, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hBC, 8'h7E, 8'h77, 8'h5C, 8'h52, 8'h62, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h51, 8'hAC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h86, 8'h5A, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h69, 8'h5E, 8'h40, 8'h5F, 8'hA6, 8'hB3, 8'hD8, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hD8, 8'hB2, 8'hA5, 8'h5F, 8'h40, 8'h5F, 8'h69, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5A, 8'h86, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h67, 8'h61, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5B, 8'h3A, 8'h67, 8'hCD, 8'hDD, 8'hEE, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hEE, 8'hDD, 8'hCB, 8'h66, 8'h3A, 8'h5C, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h61, 8'h67, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h54, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h61, 8'h5A, 8'h4D, 8'h7C, 8'hE7, 8'hF8, 8'hFB, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFB, 8'hF8, 8'hE5, 8'h7B, 8'h4D, 8'h5B, 8'h61, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h54, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h4E, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h55, 8'h5A, 8'h77, 8'h9D, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h9C, 8'h77, 8'h5B, 8'h55, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4E, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'h4F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h47, 8'h5C, 8'hAF, 8'hC5, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hC5, 8'hAF, 8'h5B, 8'h47, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4F, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'h50, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h41, 8'h62, 8'hDC, 8'hE5, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE5, 8'hDC, 8'h62, 8'h41, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h50, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'h52, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h5D, 8'h51, 8'h77, 8'hF7, 8'hF9, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF9, 8'hF7, 8'h77, 8'h50, 8'h5C, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h52, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h56, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h61, 8'h50, 8'h73, 8'h99, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h99, 8'h73, 8'h50, 8'h61, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h56, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h98, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h5E, 8'h42, 8'hA0, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC2, 8'h9F, 8'h41, 8'h5E, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'h98, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h81, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5B, 8'h3D, 8'hC5, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'hC5, 8'h3C, 8'h5B, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6D, 8'h62, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h59, 8'h51, 8'hE0, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hDF, 8'h50, 8'h59, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h62, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h60, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5D, 8'h59, 8'h7B, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'h7A, 8'h59, 8'h5D, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h60, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h55, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h54, 8'h5B, 8'hB0, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hB0, 8'h59, 8'h54, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h55, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h4C, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h50, 8'h61, 8'hDC, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hDC, 8'h60, 8'h50, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4C, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'h49, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h54, 8'h77, 8'hF7, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF7, 8'h75, 8'h54, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h49, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h4D, 8'h65, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5A, 8'h5F, 8'h99, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h97, 8'h5F, 8'h5A, 8'h67, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4D, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD7, 8'h52, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h51, 8'h70, 8'hC2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC2, 8'h70, 8'h51, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h52, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'h57, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4B, 8'h81, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'h81, 8'h4B, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h57, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h51, 8'h98, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h98, 8'h51, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAE, 8'h5C, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5D, 8'h60, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB4, 8'h61, 8'h5D, 8'h67, 8'h66, 8'h66, 8'h66, 8'h5C, 8'hAE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA3, 8'h5E, 8'h66, 8'h66, 8'h66, 8'h67, 8'h54, 8'h75, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'h75, 8'h54, 8'h67, 8'h66, 8'h66, 8'h66, 8'h5E, 8'hA3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h98, 8'h5E, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4F, 8'h8A, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFC, 8'hFB, 8'hFA, 8'hF9, 8'hF8, 8'hF8, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF8, 8'hF8, 8'hF9, 8'hFA, 8'hFB, 8'hFC, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h8A, 8'h4F, 8'h67, 8'h66, 8'h66, 8'h66, 8'h5E, 8'h99, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8F, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h65, 8'h50, 8'hA2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'hF0, 8'hEC, 8'hE7, 8'hE4, 8'hE0, 8'hDD, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDC, 8'hDC, 8'hDC, 8'hDC, 8'hDC, 8'hDC, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDD, 8'hE1, 8'hE4, 8'hE7, 8'hEC, 8'hF1, 8'hF6, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hA3, 8'h50, 8'h65, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h8F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h86, 8'h60, 8'h66, 8'h66, 8'h66, 8'h62, 8'h58, 8'hBB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hEA, 8'hDE, 8'hD4, 8'hC9, 8'hC1, 8'hB9, 8'hB2, 8'hAD, 8'hAD, 8'hAD, 8'hAE, 8'hAF, 8'hAF, 8'hAF, 8'hAF, 8'hAF, 8'hAF, 8'hAE, 8'hAD, 8'hAD, 8'hAD, 8'hB2, 8'hBA, 8'hC2, 8'hC9, 8'hD4, 8'hDF, 8'hEB, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBC, 8'h58, 8'h62, 8'h66, 8'h66, 8'h66, 8'h60, 8'h87, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h61, 8'h66, 8'h66, 8'h66, 8'h5D, 8'h64, 8'hD7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hDB, 8'hC7, 8'hB6, 8'hA5, 8'h96, 8'h89, 8'h7E, 8'h75, 8'h75, 8'h76, 8'h76, 8'h78, 8'h78, 8'h79, 8'h79, 8'h78, 8'h78, 8'h76, 8'h76, 8'h75, 8'h75, 8'h7E, 8'h8A, 8'h97, 8'hA5, 8'hB7, 8'hC8, 8'hDD, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD7, 8'h64, 8'h5D, 8'h66, 8'h66, 8'h66, 8'h61, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h77, 8'h62, 8'h66, 8'h66, 8'h66, 8'h5A, 8'h72, 8'hED, 8'hFE, 8'hFC, 8'hFA, 8'hF8, 8'hF7, 8'hF7, 8'hE6, 8'hCA, 8'hB1, 8'h9C, 8'h86, 8'h74, 8'h63, 8'h55, 8'h4A, 8'h4A, 8'h4A, 8'h4B, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4B, 8'h4A, 8'h4A, 8'h4A, 8'h55, 8'h64, 8'h75, 8'h86, 8'h9D, 8'hB3, 8'hCD, 8'hE8, 8'hF7, 8'hF7, 8'hF8, 8'hFA, 8'hFC, 8'hFE, 8'hED, 8'h72, 8'h5A, 8'h66, 8'h66, 8'h66, 8'h62, 8'h77, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h71, 8'h62, 8'h66, 8'h66, 8'h65, 8'h5A, 8'h89, 8'hFB, 8'hFB, 8'hF1, 8'hE8, 8'hE0, 8'hDB, 8'hDC, 8'hCC, 8'hB2, 8'h9A, 8'h85, 8'h70, 8'h5F, 8'h4F, 8'h41, 8'h36, 8'h37, 8'h37, 8'h38, 8'h3B, 8'h3B, 8'h3B, 8'h3B, 8'h3B, 8'h3B, 8'h38, 8'h37, 8'h37, 8'h36, 8'h41, 8'h50, 8'h60, 8'h70, 8'h86, 8'h9B, 8'hB4, 8'hCE, 8'hDC, 8'hDB, 8'hE0, 8'hE9, 8'hF1, 8'hFB, 8'hFB, 8'h89, 8'h5A, 8'h65, 8'h66, 8'h66, 8'h62, 8'h71, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6B, 8'h63, 8'h66, 8'h66, 8'h65, 8'h5D, 8'hA8, 8'hFF, 8'hF6, 8'hE0, 8'hCC, 8'hB9, 8'hAD, 8'hB0, 8'hA6, 8'h94, 8'h83, 8'h75, 8'h65, 8'h59, 8'h4E, 8'h44, 8'h3D, 8'h3D, 8'h3E, 8'h3F, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h3F, 8'h3E, 8'h3D, 8'h3D, 8'h44, 8'h4F, 8'h5A, 8'h65, 8'h75, 8'h84, 8'h96, 8'hA7, 8'hB0, 8'hAD, 8'hB9, 8'hCC, 8'hE0, 8'hF6, 8'hFF, 8'hA8, 8'h5D, 8'h65, 8'h66, 8'h66, 8'h63, 8'h6B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h66, 8'h63, 8'h66, 8'h66, 8'h63, 8'h61, 8'hCB, 8'hFF, 8'hEF, 8'hCA, 8'hA8, 8'h89, 8'h74, 8'h7A, 8'h78, 8'h71, 8'h6A, 8'h65, 8'h5F, 8'h5B, 8'h56, 8'h52, 8'h4F, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h52, 8'h52, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h4F, 8'h52, 8'h56, 8'h5B, 8'h5F, 8'h66, 8'h6B, 8'h72, 8'h79, 8'h7A, 8'h74, 8'h89, 8'hAA, 8'hCB, 8'hEF, 8'hFF, 8'hCB, 8'h61, 8'h63, 8'h66, 8'h66, 8'h63, 8'h66, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h61, 8'h64, 8'h66, 8'h66, 8'h63, 8'h66, 8'hE2, 8'hF7, 8'hE4, 8'hB5, 8'h8A, 8'h63, 8'h49, 8'h50, 8'h54, 8'h57, 8'h58, 8'h5A, 8'h5A, 8'h5C, 8'h5C, 8'h5D, 8'h5D, 8'h5E, 8'h5E, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5E, 8'h5E, 8'h5D, 8'h5D, 8'h5C, 8'h5B, 8'h5A, 8'h5A, 8'h58, 8'h57, 8'h55, 8'h50, 8'h49, 8'h63, 8'h8C, 8'hB6, 8'hE4, 8'hF7, 8'hE2, 8'h66, 8'h63, 8'h66, 8'h66, 8'h64, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5E, 8'h64, 8'h66, 8'h66, 8'h62, 8'h6F, 8'hDD, 8'hDB, 8'hCA, 8'h9D, 8'h75, 8'h4F, 8'h36, 8'h3D, 8'h44, 8'h4B, 8'h50, 8'h55, 8'h59, 8'h5E, 8'h61, 8'h63, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h63, 8'h60, 8'h5D, 8'h59, 8'h55, 8'h50, 8'h4B, 8'h44, 8'h3D, 8'h36, 8'h4F, 8'h76, 8'h9E, 8'hCA, 8'hDB, 8'hDD, 8'h6F, 8'h62, 8'h66, 8'h66, 8'h64, 8'h5E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5C, 8'h64, 8'h66, 8'h66, 8'h61, 8'h7B, 8'hBD, 8'hAD, 8'hA5, 8'h85, 8'h69, 8'h4E, 8'h3C, 8'h42, 8'h48, 8'h4E, 8'h53, 8'h58, 8'h5C, 8'h60, 8'h63, 8'h65, 8'h68, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h68, 8'h65, 8'h62, 8'h5F, 8'h5C, 8'h58, 8'h53, 8'h4E, 8'h48, 8'h42, 8'h3C, 8'h4E, 8'h6A, 8'h86, 8'hA5, 8'hAD, 8'hBD, 8'h7B, 8'h61, 8'h66, 8'h66, 8'h64, 8'h5C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5A, 8'h64, 8'h66, 8'h66, 8'h61, 8'h8A, 8'h91, 8'h74, 8'h78, 8'h6B, 8'h60, 8'h56, 8'h4F, 8'h53, 8'h56, 8'h59, 8'h5C, 8'h5E, 8'h60, 8'h63, 8'h64, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h64, 8'h63, 8'h60, 8'h5E, 8'h5C, 8'h59, 8'h56, 8'h53, 8'h4F, 8'h56, 8'h61, 8'h6B, 8'h78, 8'h74, 8'h91, 8'h8A, 8'h61, 8'h66, 8'h66, 8'h64, 8'h5A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h64, 8'h66, 8'h66, 8'h61, 8'h92, 8'h6C, 8'h49, 8'h55, 8'h57, 8'h5A, 8'h5C, 8'h5D, 8'h60, 8'h60, 8'h61, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h61, 8'h60, 8'h60, 8'h5D, 8'h5C, 8'h5A, 8'h57, 8'h55, 8'h49, 8'h6C, 8'h92, 8'h61, 8'h66, 8'h66, 8'h64, 8'h59, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h64, 8'h66, 8'h66, 8'h61, 8'h90, 8'h58, 8'h36, 8'h45, 8'h4E, 8'h58, 8'h61, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h61, 8'h58, 8'h4E, 8'h45, 8'h36, 8'h58, 8'h90, 8'h61, 8'h66, 8'h66, 8'h64, 8'h59, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5B, 8'h64, 8'h66, 8'h66, 8'h63, 8'h83, 8'h55, 8'h3C, 8'h4A, 8'h52, 8'h5B, 8'h63, 8'h68, 8'h69, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h69, 8'h68, 8'h63, 8'h5B, 8'h52, 8'h4A, 8'h3C, 8'h55, 8'h83, 8'h63, 8'h66, 8'h66, 8'h64, 8'h5B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5C, 8'h63, 8'h66, 8'h66, 8'h64, 8'h71, 8'h59, 8'h4F, 8'h56, 8'h5B, 8'h60, 8'h64, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h68, 8'h67, 8'h68, 8'h68, 8'h68, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h69, 8'h68, 8'h68, 8'h68, 8'h67, 8'h68, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h64, 8'h60, 8'h5B, 8'h56, 8'h4F, 8'h59, 8'h71, 8'h64, 8'h66, 8'h66, 8'h63, 8'h5C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5F, 8'h63, 8'h66, 8'h66, 8'h66, 8'h62, 8'h5D, 8'h5D, 8'h61, 8'h62, 8'h64, 8'h65, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h67, 8'h67, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h67, 8'h67, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h65, 8'h64, 8'h62, 8'h61, 8'h5D, 8'h5D, 8'h62, 8'h66, 8'h66, 8'h66, 8'h63, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h63, 8'h63, 8'h66, 8'h66, 8'h67, 8'h5B, 8'h60, 8'h66, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h65, 8'h64, 8'h64, 8'h62, 8'h61, 8'h61, 8'h60, 8'h60, 8'h60, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h62, 8'h64, 8'h64, 8'h65, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h66, 8'h60, 8'h5B, 8'h67, 8'h66, 8'h66, 8'h63, 8'h63, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h69, 8'h63, 8'h66, 8'h66, 8'h67, 8'h5C, 8'h62, 8'h68, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h63, 8'h60, 8'h5E, 8'h5B, 8'h59, 8'h57, 8'h55, 8'h54, 8'h53, 8'h52, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h52, 8'h53, 8'h54, 8'h55, 8'h57, 8'h59, 8'h5B, 8'h5E, 8'h60, 8'h63, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h68, 8'h62, 8'h5C, 8'h67, 8'h66, 8'h66, 8'h63, 8'h69, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6F, 8'h62, 8'h66, 8'h66, 8'h66, 8'h61, 8'h63, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h69, 8'h67, 8'h62, 8'h5C, 8'h57, 8'h52, 8'h4E, 8'h4B, 8'h48, 8'h45, 8'h43, 8'h41, 8'h41, 8'h40, 8'h3F, 8'h3F, 8'h40, 8'h41, 8'h41, 8'h43, 8'h45, 8'h48, 8'h4B, 8'h4E, 8'h52, 8'h57, 8'h5C, 8'h62, 8'h67, 8'h69, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h67, 8'h63, 8'h61, 8'h66, 8'h66, 8'h66, 8'h62, 8'h6F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h78, 8'h61, 8'h66, 8'h66, 8'h66, 8'h64, 8'h65, 8'h67, 8'h67, 8'h66, 8'h66, 8'h67, 8'h66, 8'h67, 8'h67, 8'h65, 8'h5F, 8'h59, 8'h54, 8'h4E, 8'h4B, 8'h47, 8'h43, 8'h41, 8'h3E, 8'h3B, 8'h3B, 8'h3A, 8'h38, 8'h38, 8'h3A, 8'h3B, 8'h3B, 8'h3E, 8'h41, 8'h43, 8'h47, 8'h4B, 8'h4E, 8'h54, 8'h59, 8'h5F, 8'h65, 8'h67, 8'h67, 8'h66, 8'h67, 8'h66, 8'h66, 8'h67, 8'h67, 8'h65, 8'h64, 8'h66, 8'h66, 8'h66, 8'h61, 8'h78, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h85, 8'h5E, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h66, 8'h65, 8'h63, 8'h61, 8'h60, 8'h5F, 8'h5D, 8'h5C, 8'h5A, 8'h59, 8'h57, 8'h57, 8'h55, 8'h55, 8'h54, 8'h51, 8'h4E, 8'h4E, 8'h4D, 8'h4B, 8'h4B, 8'h4D, 8'h4E, 8'h4E, 8'h51, 8'h54, 8'h55, 8'h55, 8'h56, 8'h57, 8'h59, 8'h5A, 8'h5C, 8'h5D, 8'h5F, 8'h60, 8'h61, 8'h63, 8'h65, 8'h66, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5E, 8'h85, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h96, 8'h59, 8'h67, 8'h66, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h61, 8'h5D, 8'h59, 8'h55, 8'h51, 8'h50, 8'h58, 8'h5F, 8'h66, 8'h6B, 8'h71, 8'h76, 8'h7A, 8'h7D, 8'h7B, 8'h79, 8'h78, 8'h77, 8'h76, 8'h76, 8'h77, 8'h78, 8'h79, 8'h7B, 8'h7D, 8'h7A, 8'h76, 8'h71, 8'h6B, 8'h65, 8'h5F, 8'h58, 8'h4F, 8'h51, 8'h55, 8'h59, 8'h5D, 8'h61, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h66, 8'h67, 8'h59, 8'h96, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAB, 8'h52, 8'h69, 8'h67, 8'h67, 8'h67, 8'h67, 8'h68, 8'h69, 8'h65, 8'h5E, 8'h56, 8'h4E, 8'h47, 8'h3F, 8'h40, 8'h53, 8'h65, 8'h76, 8'h86, 8'h94, 8'h9F, 8'hA9, 8'hB2, 8'hB0, 8'hAF, 8'hAF, 8'hAF, 8'hAE, 8'hAE, 8'hAF, 8'hAF, 8'hAF, 8'hB0, 8'hB2, 8'hA9, 8'h9F, 8'h93, 8'h86, 8'h76, 8'h65, 8'h53, 8'h3F, 8'h3F, 8'h47, 8'h4E, 8'h56, 8'h5E, 8'h66, 8'h69, 8'h68, 8'h67, 8'h67, 8'h67, 8'h67, 8'h69, 8'h52, 8'hAB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBD, 8'h4E, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h67, 8'h63, 8'h5B, 8'h53, 8'h4B, 8'h43, 8'h39, 8'h3A, 8'h56, 8'h70, 8'h88, 8'h9E, 8'hB2, 8'hC3, 8'hD1, 8'hDD, 8'hDC, 8'hDC, 8'hDC, 8'hDC, 8'hDB, 8'hDB, 8'hDC, 8'hDC, 8'hDC, 8'hDC, 8'hDD, 8'hD1, 8'hC3, 8'hB1, 8'h9E, 8'h87, 8'h70, 8'h56, 8'h39, 8'h39, 8'h43, 8'h4B, 8'h53, 8'h5B, 8'h64, 8'h67, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h4E, 8'hBD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'h4E, 8'h62, 8'h65, 8'h65, 8'h64, 8'h62, 8'h60, 8'h5F, 8'h5C, 8'h5B, 8'h59, 8'h57, 8'h55, 8'h4C, 8'h4D, 8'h6A, 8'h86, 8'h9F, 8'hB6, 8'hCA, 8'hDC, 8'hEB, 8'hF8, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF7, 8'hF8, 8'hEB, 8'hDC, 8'hCA, 8'hB6, 8'h9E, 8'h86, 8'h6A, 8'h4C, 8'h4C, 8'h55, 8'h57, 8'h59, 8'h5B, 8'h5D, 8'h5F, 8'h61, 8'h62, 8'h64, 8'h65, 8'h65, 8'h62, 8'h4E, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'h52, 8'h58, 8'h61, 8'h63, 8'h60, 8'h5B, 8'h56, 8'h51, 8'h51, 8'h5D, 8'h68, 8'h72, 8'h7B, 8'h77, 8'h78, 8'h8F, 8'hA5, 8'hB9, 8'hCB, 8'hDB, 8'hE9, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hE9, 8'hDB, 8'hCB, 8'hB8, 8'hA5, 8'h8F, 8'h77, 8'h77, 8'h7B, 8'h72, 8'h68, 8'h5D, 8'h51, 8'h51, 8'h56, 8'h5B, 8'h60, 8'h63, 8'h61, 8'h58, 8'h52, 8'hDC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h59, 8'h4B, 8'h5E, 8'h61, 8'h5B, 8'h51, 8'h48, 8'h3F, 8'h43, 8'h60, 8'h7B, 8'h95, 8'hAD, 8'hAE, 8'hAF, 8'hBC, 8'hC9, 8'hD5, 8'hE0, 8'hEA, 8'hF2, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF2, 8'hE9, 8'hE0, 8'hD5, 8'hC9, 8'hBC, 8'hAE, 8'hAE, 8'hAD, 8'h95, 8'h7B, 8'h60, 8'h43, 8'h3F, 8'h4A, 8'h51, 8'h5B, 8'h61, 8'h5E, 8'h4B, 8'h59, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h64, 8'h46, 8'h5B, 8'h5E, 8'h58, 8'h4E, 8'h44, 8'h39, 8'h3F, 8'h68, 8'h8F, 8'hB4, 8'hD6, 8'hDB, 8'hDC, 8'hE2, 8'hE7, 8'hED, 8'hF1, 8'hF6, 8'hF9, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF9, 8'hF5, 8'hF1, 8'hEC, 8'hE7, 8'hE2, 8'hDB, 8'hDB, 8'hD6, 8'hB4, 8'h8F, 8'h68, 8'h3F, 8'h39, 8'h46, 8'h4E, 8'h58, 8'h5E, 8'h5B, 8'h46, 8'h64, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h7B, 8'h51, 8'h5A, 8'h5B, 8'h5A, 8'h57, 8'h54, 8'h4C, 8'h53, 8'h7E, 8'hA6, 8'hCC, 8'hF0, 8'hF7, 8'hF7, 8'hF9, 8'hFA, 8'hFB, 8'hFC, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFD, 8'hFC, 8'hFB, 8'hFA, 8'hF9, 8'hF7, 8'hF7, 8'hF0, 8'hCC, 8'hA6, 8'h7E, 8'h52, 8'h4C, 8'h56, 8'h57, 8'h5A, 8'h5B, 8'h5A, 8'h51, 8'h7B, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9C, 8'h6B, 8'h5C, 8'h59, 8'h61, 8'h6D, 8'h78, 8'h77, 8'h7C, 8'h9E, 8'hBE, 8'hDC, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hDC, 8'hBE, 8'h9E, 8'h7C, 8'h77, 8'h79, 8'h6D, 8'h61, 8'h59, 8'h5C, 8'h6B, 8'h9C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h8C, 8'h5F, 8'h55, 8'h6A, 8'h88, 8'hA6, 8'hAE, 8'hB2, 8'hC6, 8'hD9, 8'hEB, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hEB, 8'hD9, 8'hC6, 8'hB1, 8'hAE, 8'hA6, 8'h88, 8'h6A, 8'h55, 8'h5F, 8'h8C, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hAB, 8'h67, 8'h59, 8'h76, 8'hA2, 8'hCC, 8'hDB, 8'hDD, 8'hE6, 8'hEE, 8'hF6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF6, 8'hEE, 8'hE6, 8'hDD, 8'hDB, 8'hCC, 8'hA2, 8'h76, 8'h59, 8'h67, 8'hAB, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC4, 8'h7C, 8'h6E, 8'h8C, 8'hBA, 8'hE6, 8'hF7, 8'hF8, 8'hF9, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hF9, 8'hF7, 8'hF7, 8'hE5, 8'hBA, 8'h8C, 8'h6E, 8'h7C, 8'hC4, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h9D, 8'h92, 8'hAA, 8'hCE, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hCE, 8'hAA, 8'h92, 8'h9D, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hC5, 8'hBE, 8'hCC, 8'hE2, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hE2, 8'hCC, 8'hBE, 8'hC5, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE5, 8'hE2, 8'hE9, 8'hF2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF2, 8'hE9, 8'hE2, 8'hE5, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF9, 8'hF9, 8'hFA, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hFA, 8'hF9, 8'hF9, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hE8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hE8, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF7, 8'hE1, 8'hDA, 8'hF7, 8'hF8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF8, 8'hF7, 8'hDA, 8'hE1, 8'hF7, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'hDA, 8'hC7, 8'hC1, 8'hDC, 8'hDD, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hDD, 8'hDC, 8'hC1, 8'hC7, 8'hDA, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hAC, 8'hA3, 8'h9E, 8'hB0, 8'hB2, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hB2, 8'hB0, 8'h9E, 8'hA3, 8'hAC, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA0, 8'h73, 8'h77, 8'h75, 8'h7B, 8'h7C, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h7C, 8'h7B, 8'h75, 8'h77, 8'h73, 8'hA0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h7F, 8'h47, 8'h56, 8'h55, 8'h51, 8'h53, 8'hE6, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hE6, 8'h53, 8'h51, 8'h55, 8'h56, 8'h47, 8'h80, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h69, 8'h34, 8'h46, 8'h47, 8'h3F, 8'h3F, 8'hCA, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hCA, 8'h3F, 8'h3F, 8'h47, 8'h46, 8'h34, 8'h6A, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h60, 8'h3C, 8'h4A, 8'h4B, 8'h44, 8'h43, 8'hA0, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hA0, 8'h43, 8'h44, 8'h4B, 8'h4A, 8'h3C, 8'h60, 8'hB7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h86, 8'h5A, 8'h4E, 8'h57, 8'h57, 8'h53, 8'h51, 8'h6F, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h6F, 8'h51, 8'h53, 8'h57, 8'h57, 8'h4E, 8'h5B, 8'h86, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h5E, 8'h57, 8'h5E, 8'h61, 8'h61, 8'h60, 8'h5C, 8'h48, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h48, 8'h5C, 8'h60, 8'h61, 8'h61, 8'h5E, 8'h57, 8'h5E, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'h49, 8'h57, 8'h67, 8'h67, 8'h67, 8'h67, 8'h63, 8'h38, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'h38, 8'h63, 8'h67, 8'h67, 8'h67, 8'h67, 8'h57, 8'h49, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE1, 8'h46, 8'h5B, 8'h69, 8'h68, 8'h68, 8'h69, 8'h65, 8'h3E, 8'hAB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAB, 8'h3E, 8'h65, 8'h69, 8'h68, 8'h68, 8'h69, 8'h5B, 8'h46, 8'hE1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'h4C, 8'h60, 8'h67, 8'h67, 8'h67, 8'h67, 8'h66, 8'h4F, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h80, 8'h4F, 8'h66, 8'h67, 8'h67, 8'h67, 8'h67, 8'h60, 8'h4C, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB9, 8'h51, 8'h64, 8'h67, 8'h66, 8'h66, 8'h67, 8'h66, 8'h5C, 8'h5E, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h5E, 8'h5C, 8'h66, 8'h67, 8'h66, 8'h66, 8'h67, 8'h64, 8'h51, 8'hB9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA5, 8'h56, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h4A, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'h4A, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h56, 8'hA5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h5A, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h48, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'h48, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5A, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h5D, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4B, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'h4B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5D, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6E, 8'h61, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4F, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'h4F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h61, 8'h6E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h61, 8'h63, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h52, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h52, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h63, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h55, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'h55, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h59, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h58, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'h58, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4E, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5A, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h5A, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4C, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4D, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5C, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB4, 8'h5C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB4, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h4F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h51, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h51, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h53, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h52, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h52, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h50, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5B, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h5B, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h50, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4D, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5C, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h5C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4C, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5C, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB4, 8'h5C, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4E, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5A, 8'hB9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB9, 8'h5A, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h4E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h53, 8'h65, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h59, 8'hC1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC1, 8'h59, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h65, 8'h52, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h58, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h56, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'h56, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h57, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h60, 8'h64, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h54, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h54, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h64, 8'h5E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h62, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h50, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'h50, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h62, 8'h6A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7B, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h4C, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'h4C, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h5B, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h68, 8'h46, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'h46, 8'h68, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h5B, 8'h8C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9F, 8'h57, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h48, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h48, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h66, 8'h57, 8'h9E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h51, 8'h65, 8'h67, 8'h66, 8'h66, 8'h66, 8'h66, 8'h5F, 8'h5A, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h5A, 8'h5F, 8'h66, 8'h66, 8'h66, 8'h66, 8'h67, 8'h65, 8'h51, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'h4A, 8'h61, 8'h68, 8'h67, 8'h67, 8'h67, 8'h66, 8'h52, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h52, 8'h66, 8'h67, 8'h67, 8'h67, 8'h68, 8'h61, 8'h4A, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h42, 8'h5E, 8'h69, 8'h68, 8'h68, 8'h68, 8'h67, 8'h41, 8'hA3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA3, 8'h41, 8'h67, 8'h68, 8'h68, 8'h68, 8'h69, 8'h5E, 8'h42, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h42, 8'h5A, 8'h68, 8'h67, 8'h67, 8'h67, 8'h65, 8'h3B, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h3B, 8'h65, 8'h67, 8'h67, 8'h67, 8'h68, 8'h5A, 8'h42, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h58, 8'h58, 8'h60, 8'h62, 8'h62, 8'h60, 8'h5C, 8'h49, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h49, 8'h5C, 8'h60, 8'h62, 8'h62, 8'h60, 8'h58, 8'h58, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h81, 8'h57, 8'h51, 8'h58, 8'h59, 8'h55, 8'h4F, 8'h6B, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'h6B, 8'h4F, 8'h55, 8'h59, 8'h58, 8'h51, 8'h57, 8'h81, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB4, 8'h57, 8'h40, 8'h4D, 8'h4D, 8'h47, 8'h3E, 8'h97, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'h97, 8'h3E, 8'h47, 8'h4D, 8'h4D, 8'h40, 8'h57, 8'hB4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h5C, 8'h39, 8'h49, 8'h49, 8'h43, 8'h38, 8'hBD, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hBD, 8'h38, 8'h43, 8'h49, 8'h49, 8'h39, 8'h5C, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h72, 8'h4C, 8'h56, 8'h56, 8'h53, 8'h4C, 8'hD8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hD8, 8'h4C, 8'h53, 8'h56, 8'h56, 8'h4C, 8'h72, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h77, 8'h74, 8'h72, 8'h78, 8'h77, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h77, 8'h78, 8'h72, 8'h74, 8'h77, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC0, 8'hAE, 8'h9A, 8'h96, 8'hA8, 8'hAE, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hAE, 8'hA8, 8'h96, 8'h9A, 8'hAE, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hDB, 8'hBB, 8'hB6, 8'hCF, 8'hDB, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hDB, 8'hCF, 8'hB6, 8'hBB, 8'hDB, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF7, 8'hD4, 8'hCE, 8'hE9, 8'hF7, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF7, 8'hE9, 8'hCE, 8'hD4, 8'hF7, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hDE, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDE, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hEC, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hEC, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hF6, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF6, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF}; 
reg	[7:0]	pattern_data_B1 [0:39999] = '{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF9, 8'hF8, 8'hF8, 8'hF9, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hF2, 8'hF0, 8'hF0, 8'hF2, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hE9, 8'hE5, 8'hE5, 8'hE9, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hF9, 8'hF7, 8'hF6, 8'hF6, 8'hF6, 8'hE7, 8'hDB, 8'hD6, 8'hD6, 8'hDB, 8'hE7, 8'hF6, 8'hF6, 8'hF6, 8'hF7, 8'hF9, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hEB, 8'hE1, 8'hD9, 8'hD5, 8'hD6, 8'hD8, 8'hC9, 8'hBD, 8'hB8, 8'hB8, 8'hBD, 8'hC9, 8'hD8, 8'hD6, 8'hD5, 8'hD9, 8'hE1, 8'hEB, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hD1, 8'hBC, 8'hA8, 8'hA0, 8'hA3, 8'hA6, 8'h9B, 8'h93, 8'h8F, 8'h8F, 8'h93, 8'h9B, 8'hA6, 8'hA3, 8'hA0, 8'hA8, 8'hBC, 8'hD1, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB2, 8'h8D, 8'h6D, 8'h5F, 8'h63, 8'h68, 8'h64, 8'h60, 8'h5F, 8'h5F, 8'h60, 8'h64, 8'h68, 8'h63, 8'h5F, 8'h6D, 8'h8D, 8'hB2, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF9, 8'hF6, 8'hF6, 8'hC8, 8'h95, 8'h67, 8'h3E, 8'h2D, 8'h32, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h32, 8'h2D, 8'h3E, 8'h67, 8'h95, 8'hC9, 8'hF6, 8'hF6, 8'hF9, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hE5, 8'hD7, 8'hD7, 8'hAB, 8'h7B, 8'h4E, 8'h27, 8'h16, 8'h1C, 8'h22, 8'h25, 8'h27, 8'h28, 8'h28, 8'h27, 8'h25, 8'h22, 8'h1C, 8'h16, 8'h27, 8'h4E, 8'h7B, 8'hAC, 8'hD6, 8'hD7, 8'hE6, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hC5, 8'hA4, 8'hA3, 8'h86, 8'h64, 8'h45, 8'h2A, 8'h1E, 8'h23, 8'h28, 8'h2A, 8'h2C, 8'h2D, 8'h2D, 8'h2C, 8'h2A, 8'h28, 8'h23, 8'h1E, 8'h2A, 8'h45, 8'h64, 8'h87, 8'hA3, 8'hA4, 8'hC5, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h9C, 8'h65, 8'h64, 8'h5B, 8'h4F, 8'h42, 8'h37, 8'h33, 8'h35, 8'h38, 8'h3A, 8'h3B, 8'h3B, 8'h3B, 8'h3B, 8'h3A, 8'h38, 8'h35, 8'h33, 8'h37, 8'h42, 8'h4F, 8'h5C, 8'h63, 8'h65, 8'h9E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF8, 8'hF6, 8'hC8, 8'h7A, 8'h35, 8'h33, 8'h3A, 8'h3E, 8'h40, 8'h42, 8'h44, 8'h45, 8'h46, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h46, 8'h45, 8'h44, 8'h42, 8'h40, 8'h3E, 8'h3B, 8'h32, 8'h35, 8'h7C, 8'hC9, 8'hF6, 8'hF8, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hE1, 8'hD5, 8'hAB, 8'h61, 8'h1E, 8'h1D, 8'h2B, 8'h37, 8'h40, 8'h49, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h49, 8'h40, 8'h37, 8'h2B, 8'h1C, 8'h1E, 8'h62, 8'hAC, 8'hD5, 8'hE1, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hBB, 8'hA0, 8'h86, 8'h52, 8'h23, 8'h24, 8'h30, 8'h3B, 8'h43, 8'h4C, 8'h50, 8'h50, 8'h50, 8'h50, 8'h4F, 8'h4F, 8'h4F, 8'h4F, 8'h50, 8'h50, 8'h50, 8'h50, 8'h4C, 8'h43, 8'h3B, 8'h30, 8'h23, 8'h23, 8'h53, 8'h87, 8'hA0, 8'hBB, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h8C, 8'h5F, 8'h5B, 8'h47, 8'h34, 8'h36, 8'h3D, 8'h43, 8'h48, 8'h4C, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4C, 8'h48, 8'h43, 8'h3D, 8'h36, 8'h34, 8'h48, 8'h5C, 8'h5F, 8'h8D, 8'hDC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF6, 8'hC9, 8'h65, 8'h2D, 8'h3A, 8'h3F, 8'h42, 8'h46, 8'h48, 8'h4A, 8'h4B, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4B, 8'h4A, 8'h48, 8'h46, 8'h42, 8'h3F, 8'h3B, 8'h2D, 8'h66, 8'hCA, 8'hF6, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hD6, 8'hAC, 8'h4C, 8'h16, 8'h2B, 8'h3C, 8'h4B, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4B, 8'h3C, 8'h2B, 8'h16, 8'h4E, 8'hAD, 8'hD6, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hA1, 8'h87, 8'h43, 8'h1E, 8'h30, 8'h40, 8'h4D, 8'h50, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4F, 8'h50, 8'h4D, 8'h40, 8'h30, 8'h1E, 8'h45, 8'h87, 8'hA1, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h60, 8'h5C, 8'h41, 8'h33, 8'h3D, 8'h45, 8'h4D, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4F, 8'h4D, 8'h45, 8'h3D, 8'h33, 8'h41, 8'h5C, 8'h60, 8'hAE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF6, 8'h8F, 8'h2E, 8'h3B, 8'h3F, 8'h44, 8'h48, 8'h4A, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h4A, 8'h48, 8'h44, 8'h40, 8'h3A, 8'h2E, 8'h90, 8'hF6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'hD5, 8'h74, 8'h18, 8'h2B, 8'h40, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h40, 8'h2B, 8'h18, 8'h76, 8'hD5, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC1, 8'hA0, 8'h60, 8'h1F, 8'h30, 8'h43, 8'h50, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h50, 8'h43, 8'h2F, 8'h1F, 8'h61, 8'hA0, 8'hC2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h97, 8'h5F, 8'h4C, 8'h33, 8'h3D, 8'h48, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h48, 8'h3D, 8'h33, 8'h4D, 8'h5F, 8'h98, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF6, 8'h73, 8'h2D, 8'h3E, 8'h43, 8'h48, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h47, 8'h43, 8'h3E, 8'h2D, 8'h75, 8'hF6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hD5, 8'h5A, 8'h16, 8'h38, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h38, 8'h16, 8'h5B, 8'hD5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'hA0, 8'h4D, 8'h1E, 8'h3C, 8'h4F, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h4F, 8'h3C, 8'h1E, 8'h4E, 8'hA0, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9B, 8'h60, 8'h45, 8'h33, 8'h43, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h43, 8'h33, 8'h46, 8'h60, 8'h9C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'h79, 8'h2D, 8'h3F, 8'h44, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h44, 8'h3F, 8'h2D, 8'h79, 8'hF6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hD5, 8'h5F, 8'h17, 8'h3E, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h3E, 8'h17, 8'h60, 8'hD5, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'hA0, 8'h50, 8'h1F, 8'h41, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h41, 8'h1F, 8'h51, 8'hA0, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBE, 8'h5F, 8'h46, 8'h33, 8'h46, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h46, 8'h33, 8'h46, 8'h5F, 8'hBE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hA4, 8'h2D, 8'h3E, 8'h44, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h44, 8'h3E, 8'h2D, 8'hA5, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'h88, 8'h16, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'h16, 8'h89, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA9, 8'h6D, 8'h1E, 8'h3F, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h3F, 8'h1E, 8'h6E, 8'hA9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6F, 8'h50, 8'h33, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h33, 8'h50, 8'h6F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'h40, 8'h3A, 8'h44, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h44, 8'h3A, 8'h40, 8'hF6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hD6, 8'h29, 8'h31, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h31, 8'h29, 8'hD6, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hA1, 8'h2B, 8'h36, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h36, 8'h2B, 8'hA1, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB8, 8'h60, 8'h37, 8'h40, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h40, 8'h37, 8'h60, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h9D, 8'h2E, 8'h41, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h41, 8'h2E, 8'h9D, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'h81, 8'h18, 8'h48, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h48, 8'h18, 8'h81, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h67, 8'h1F, 8'h4A, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h4A, 8'h1F, 8'h67, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7E, 8'h4D, 8'h34, 8'h4C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4C, 8'h34, 8'h4B, 8'h7E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h54, 8'h39, 8'h44, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h44, 8'h37, 8'h54, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h3C, 8'h31, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h2F, 8'h3C, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA3, 8'h38, 8'h36, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h34, 8'h37, 8'hA3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h63, 8'h3B, 8'h40, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h40, 8'h3A, 8'h63, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF6, 8'h32, 8'h3F, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h3D, 8'h32, 8'hF6, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hD5, 8'h1B, 8'h43, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h41, 8'h1B, 8'hD5, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hA0, 8'h21, 8'h46, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h45, 8'h21, 8'hA0, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'h5F, 8'h32, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4E, 8'h4F, 8'h4F, 8'h4F, 8'h4F, 8'h4E, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h48, 8'h32, 8'h5F, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hDA, 8'h2D, 8'h41, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4C, 8'h4F, 8'h4F, 8'h50, 8'h50, 8'h4F, 8'h4F, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h41, 8'h2D, 8'hDA, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBB, 8'h17, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h51, 8'h51, 8'h50, 8'h50, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h17, 8'hBB, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h8D, 8'h1F, 8'h4C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4F, 8'h52, 8'h55, 8'h57, 8'h57, 8'h54, 8'h51, 8'h50, 8'h50, 8'h51, 8'h54, 8'h57, 8'h57, 8'h55, 8'h52, 8'h4F, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4C, 8'h1F, 8'h8D, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h57, 8'h33, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h52, 8'h58, 8'h5D, 8'h60, 8'h5E, 8'h58, 8'h53, 8'h50, 8'h50, 8'h53, 8'h58, 8'h60, 8'h60, 8'h5C, 8'h58, 8'h52, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h33, 8'h57, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC2, 8'h2D, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h53, 8'h59, 8'h5F, 8'h63, 8'h61, 8'h57, 8'h50, 8'h4C, 8'h4C, 8'h50, 8'h57, 8'h63, 8'h63, 8'h5E, 8'h59, 8'h53, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h2D, 8'hC1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hA4, 8'h1C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h50, 8'h51, 8'h54, 8'h55, 8'h59, 8'h58, 8'h4D, 8'h46, 8'h42, 8'h42, 8'h46, 8'h4D, 8'h59, 8'h59, 8'h55, 8'h54, 8'h51, 8'h50, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h1C, 8'hA2, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE2, 8'h7D, 8'h24, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h51, 8'h55, 8'h55, 8'h4D, 8'h47, 8'h41, 8'h44, 8'h43, 8'h3A, 8'h35, 8'h32, 8'h32, 8'h35, 8'h3A, 8'h44, 8'h44, 8'h41, 8'h47, 8'h4D, 8'h55, 8'h55, 8'h51, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h24, 8'h7C, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'h51, 8'h36, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h54, 8'h5D, 8'h5D, 8'h48, 8'h36, 8'h27, 8'h28, 8'h27, 8'h23, 8'h1F, 8'h1D, 8'h1D, 8'h1F, 8'h23, 8'h28, 8'h28, 8'h28, 8'h36, 8'h48, 8'h5D, 8'h5D, 8'h54, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h36, 8'h50, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hB9, 8'h2F, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h55, 8'h5F, 8'h5F, 8'h41, 8'h28, 8'h12, 8'h12, 8'h11, 8'h0F, 8'h0E, 8'h0D, 8'h0D, 8'h0E, 8'h0F, 8'h12, 8'h12, 8'h13, 8'h28, 8'h41, 8'h5F, 8'h5F, 8'h55, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h2F, 8'hB9, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h9B, 8'h21, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h50, 8'h52, 8'h55, 8'h55, 8'h36, 8'h1B, 8'h05, 8'h04, 8'h04, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h04, 8'h04, 8'h06, 8'h1B, 8'h36, 8'h55, 8'h55, 8'h52, 8'h50, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h21, 8'h9B, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h76, 8'h28, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h54, 8'h55, 8'h4A, 8'h41, 8'h41, 8'h28, 8'h13, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h13, 8'h28, 8'h41, 8'h41, 8'h4A, 8'h55, 8'h54, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h28, 8'h76, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h4E, 8'h39, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4E, 8'h5A, 8'h5D, 8'h40, 8'h26, 8'h26, 8'h18, 8'h0B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h0B, 8'h18, 8'h26, 8'h26, 8'h40, 8'h5D, 8'h5A, 8'h4E, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h39, 8'h4E, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC2, 8'h2E, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4F, 8'h5C, 8'h5F, 8'h36, 8'h11, 8'h11, 8'h0A, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h0A, 8'h11, 8'h11, 8'h36, 8'h5F, 8'h5C, 8'h4F, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h2E, 8'hC2, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hA3, 8'h22, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h50, 8'h55, 8'h55, 8'h2A, 8'h04, 8'h04, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h04, 8'h04, 8'h2A, 8'h55, 8'h55, 8'h50, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h22, 8'hA3, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'h7C, 8'h29, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h55, 8'h52, 8'h44, 8'h41, 8'h1F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1F, 8'h41, 8'h44, 8'h52, 8'h55, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h29, 8'h7C, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'h4F, 8'h3A, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4E, 8'h5D, 8'h55, 8'h2F, 8'h26, 8'h12, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h12, 8'h26, 8'h2F, 8'h55, 8'h5D, 8'h4E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h3A, 8'h4F, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h2C, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4F, 8'h5F, 8'h53, 8'h1D, 8'h11, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h11, 8'h1D, 8'h53, 8'h5F, 8'h4F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h2C, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h1F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h51, 8'h56, 8'h49, 8'h10, 8'h04, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h04, 8'h10, 8'h49, 8'h56, 8'h51, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h1F, 8'hBB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h27, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h53, 8'h54, 8'h44, 8'h37, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h37, 8'h44, 8'h54, 8'h53, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h27, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h57, 8'h38, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4B, 8'h58, 8'h58, 8'h2B, 8'h21, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h21, 8'h2B, 8'h58, 8'h58, 8'h4B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h38, 8'h57, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h2D, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h5A, 8'h57, 8'h17, 8'h0E, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h0E, 8'h17, 8'h57, 8'h5A, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h2D, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'h1B, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h55, 8'h4D, 8'h0A, 8'h03, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h03, 8'h0A, 8'h4D, 8'h55, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h1B, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA6, 8'h22, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4E, 8'h57, 8'h48, 8'h3A, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h3A, 8'h48, 8'h57, 8'h4E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h22, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h35, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4F, 8'h60, 8'h37, 8'h23, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h23, 8'h37, 8'h60, 8'h4F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h35, 8'h68, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h38, 8'h43, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h50, 8'h63, 8'h29, 8'h0F, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h0F, 8'h29, 8'h63, 8'h50, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h43, 8'h38, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h21, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h52, 8'h5A, 8'h1C, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h1C, 8'h5A, 8'h52, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h21, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h23, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h51, 8'h53, 8'h44, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h44, 8'h53, 8'h51, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h24, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h80, 8'h32, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h55, 8'h54, 8'h29, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h29, 8'h54, 8'h55, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h33, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h55, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h57, 8'h52, 8'h12, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h12, 8'h52, 8'h57, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'h55, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'h3B, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h54, 8'h48, 8'h04, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h04, 8'h48, 8'h54, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h3B, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h34, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h54, 8'h4C, 8'h36, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h36, 8'h4C, 8'h54, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h34, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h34, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h5C, 8'h42, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h42, 8'h5C, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h35, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9F, 8'h35, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5F, 8'h38, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h38, 8'h5F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h36, 8'h9F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h81, 8'h38, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h58, 8'h2C, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h2C, 8'h58, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h39, 8'h81, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h63, 8'h3E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h49, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h49, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h3F, 8'h63, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h44, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h5E, 8'h34, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h34, 8'h5E, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h44, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'h2C, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h61, 8'h23, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h23, 8'h61, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h2C, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h24, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h59, 8'h16, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h16, 8'h59, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h24, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h2B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h46, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h46, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h2B, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h39, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h5D, 8'h2D, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h2D, 8'h5D, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h39, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h48, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h61, 8'h19, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h19, 8'h61, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h48, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'h2F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h59, 8'h0B, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h0B, 8'h59, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h2F, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h2C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h54, 8'h46, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h46, 8'h54, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h2C, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC0, 8'h32, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5C, 8'h2F, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h2F, 8'h5C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h32, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA7, 8'h38, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5F, 8'h1B, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h1B, 8'h5F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h38, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h89, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h59, 8'h0D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0D, 8'h59, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'h88, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6A, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h4B, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h4B, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h69, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h48, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h57, 8'h39, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h38, 8'h57, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h48, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h2E, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5A, 8'h29, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h28, 8'h5A, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h2E, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h24, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h58, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1B, 8'h58, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h24, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'h29, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h52, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h12, 8'h52, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h29, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9E, 8'h35, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h50, 8'h4A, 8'h0B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0B, 8'h4A, 8'h50, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h35, 8'h9E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7C, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h51, 8'h41, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h41, 8'h51, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'h7C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5F, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h54, 8'h35, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h35, 8'h54, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h46, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4B, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h27, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h4B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3A, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h17, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h17, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h2D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h58, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h06, 8'h08, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h08, 8'h06, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h58, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h2D, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'h29, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h4D, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0D, 8'h1A, 8'h25, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h25, 8'h1A, 8'h0D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h4D, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h29, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1D, 8'h3C, 8'h55, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h55, 8'h3B, 8'h1D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9D, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h23, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h65, 8'h8F, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'h8F, 8'h64, 8'h31, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h23, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'h9D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5C, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h08, 8'h09, 8'h09, 8'h48, 8'h8A, 8'hC0, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hC0, 8'h88, 8'h48, 8'h09, 8'h09, 8'h08, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h5C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h7A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5E, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h5A, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0D, 8'h25, 8'h2A, 8'h2A, 8'h68, 8'hAB, 8'hE0, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hE0, 8'hA9, 8'h68, 8'h2A, 8'h2A, 8'h25, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h5A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h5E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4B, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1D, 8'h53, 8'h5F, 8'h5F, 8'h90, 8'hC4, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC3, 8'h90, 8'h5F, 8'h5F, 8'h53, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h4B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3A, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h8D, 8'hA0, 8'hA0, 8'hBD, 8'hDC, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hDB, 8'hBD, 8'hA0, 8'hA0, 8'h8D, 8'h2F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4A, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h2E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h09, 8'h47, 8'hBC, 8'hD5, 8'hD5, 8'hE2, 8'hF0, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hEF, 8'hE2, 8'hD5, 8'hD5, 8'hBC, 8'h45, 8'h09, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h40, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h2E, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h2A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h34, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h23, 8'h2A, 8'h67, 8'hDD, 8'hF6, 8'hF6, 8'hF9, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hF9, 8'hF6, 8'hF6, 8'hDD, 8'h66, 8'h2A, 8'h23, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h34, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2A, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h26, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4F, 8'h5F, 8'h8F, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'h8E, 8'h5F, 8'h4F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h26, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h38, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h16, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h86, 8'hA0, 8'hBD, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hBC, 8'hA0, 8'h85, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h16, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h38, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h40, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5B, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h09, 8'hB4, 8'hD5, 8'hE2, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hE2, 8'hD5, 8'hB3, 8'h09, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h5B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h40, 8'h95, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h79, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h58, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2A, 8'h2A, 8'hD4, 8'hF6, 8'hF9, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF9, 8'hF6, 8'hD3, 8'h2A, 8'h2A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h58, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h79, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h60, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h5F, 8'h5F, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'h5F, 8'h5F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h60, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h47, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hA0, 8'hA0, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hA0, 8'hA0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h47, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h09, 8'hD5, 8'hD5, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD5, 8'hD5, 8'h09, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h2B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h30, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h2A, 8'hF6, 8'hF6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF6, 8'hF6, 8'h2A, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2B, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h2D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4A, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5F, 8'h49, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2D, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h34, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h55, 8'h16, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7C, 8'hA0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA0, 8'h7C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h16, 8'h55, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h34, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'h3A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h0B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'hA8, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hA7, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0B, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3A, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB0, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h57, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2A, 8'hC8, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hC7, 8'h2A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h57, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hAF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9A, 8'h41, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h55, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h5F, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h5F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h55, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h41, 8'h99, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h81, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hA0, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hA0, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h09, 8'hD5, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hD5, 8'h09, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h46, 8'h6B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h58, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h2A, 8'hF6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF6, 8'h2A, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h57, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h49, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h43, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5F, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h43, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3B, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hA0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA0, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h30, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h31, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h32, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'h32, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h30, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'h2C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h2A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0B, 8'h53, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h53, 8'h0B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2A, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2C, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1A, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h1A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'h36, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h1E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2B, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h2B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1E, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h36, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC0, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h19, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h40, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hFA, 8'hF8, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF8, 8'hFA, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h40, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h19, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAF, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h14, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h61, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hEF, 8'hE6, 8'hDF, 8'hD8, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD8, 8'hDF, 8'hE6, 8'hF0, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h61, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h14, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hAE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9F, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h8A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hDB, 8'hC7, 8'hB6, 8'hA6, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA6, 8'hB6, 8'hC7, 8'hDC, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8A, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h9F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8F, 8'h43, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0D, 8'hBA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'hC2, 8'hA1, 8'h84, 8'h68, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h68, 8'h85, 8'hA1, 8'hC4, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h0D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h43, 8'h8F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h19, 8'hE1, 8'hFD, 8'hFA, 8'hF7, 8'hF6, 8'hF6, 8'hF6, 8'hD6, 8'hA8, 8'h7E, 8'h59, 8'h36, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h2A, 8'h36, 8'h5A, 8'h7E, 8'hAB, 8'hD6, 8'hF6, 8'hF6, 8'hF6, 8'hF7, 8'hFA, 8'hFD, 8'hE1, 8'h19, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6E, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'hF8, 8'hF7, 8'hE8, 8'hD9, 8'hD5, 8'hD5, 8'hD5, 8'hB5, 8'h88, 8'h5D, 8'h38, 8'h15, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h09, 8'h15, 8'h39, 8'h5D, 8'h8A, 8'hB5, 8'hD5, 8'hD5, 8'hD5, 8'hD9, 8'hE8, 8'hF8, 8'hF8, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h6E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5D, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h6B, 8'hFF, 8'hEE, 8'hCA, 8'hA9, 8'hA0, 8'hA0, 8'hA0, 8'h87, 8'h63, 8'h42, 8'h25, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h26, 8'h42, 8'h65, 8'h87, 8'hA0, 8'hA0, 8'hA0, 8'hA9, 8'hCA, 8'hEE, 8'hFF, 8'h6B, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h5D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4C, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hA8, 8'hFF, 8'hE2, 8'hA6, 8'h6E, 8'h5F, 8'h5F, 8'h5F, 8'h50, 8'h3B, 8'h27, 8'h16, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h16, 8'h27, 8'h3C, 8'h50, 8'h5F, 8'h5F, 8'h5F, 8'h6E, 8'hA6, 8'hE3, 8'hFF, 8'hA8, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h4B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h3D, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'hCF, 8'hF6, 8'hD1, 8'h84, 8'h3D, 8'h2A, 8'h2A, 8'h2A, 8'h23, 8'h1A, 8'h11, 8'h0A, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h0A, 8'h11, 8'h1A, 8'h23, 8'h2A, 8'h2A, 8'h2A, 8'h3D, 8'h84, 8'hD2, 8'hF6, 8'hCF, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h3C, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h35, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'hCD, 8'hD5, 8'hB0, 8'h64, 8'h1C, 8'h09, 8'h09, 8'h09, 8'h08, 8'h06, 8'h04, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h04, 8'h06, 8'h08, 8'h09, 8'h09, 8'h09, 8'h1C, 8'h64, 8'hB1, 8'hD5, 8'hCD, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h34, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'h33, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h23, 8'hA0, 8'hA0, 8'h83, 8'h47, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h47, 8'h84, 8'hA0, 8'hA0, 8'h23, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h32, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h35, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'h5F, 8'h5F, 8'h4E, 8'h2A, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h2A, 8'h4E, 8'h5F, 8'h5F, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h36, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4A, 8'h2A, 8'h2A, 8'h22, 8'h13, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h13, 8'h22, 8'h2A, 8'h2A, 8'h4A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h35, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'h37, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4A, 8'h09, 8'h09, 8'h08, 8'h04, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h04, 8'h08, 8'h09, 8'h09, 8'h4A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h37, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h23, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h23, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBF, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hBE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA7, 8'h41, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h41, 8'hA7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9C, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h06, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h9C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h43, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h01, 8'h02, 8'h02, 8'h02, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h03, 8'h02, 8'h02, 8'h02, 8'h01, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h43, 8'h92, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h87, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h05, 8'h07, 8'h09, 8'h0B, 8'h0C, 8'h0D, 8'h0E, 8'h0F, 8'h0F, 8'h0F, 8'h0F, 8'h0F, 8'h0F, 8'h0E, 8'h0D, 8'h0C, 8'h0B, 8'h09, 8'h07, 8'h05, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0F, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h88, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7E, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h17, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h07, 8'h0C, 8'h11, 8'h15, 8'h19, 8'h1C, 8'h1E, 8'h20, 8'h21, 8'h23, 8'h23, 8'h23, 8'h23, 8'h21, 8'h20, 8'h1E, 8'h1C, 8'h19, 8'h15, 8'h11, 8'h0C, 8'h07, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h17, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h0B, 8'h14, 8'h1C, 8'h23, 8'h2A, 8'h2E, 8'h33, 8'h37, 8'h38, 8'h3A, 8'h3B, 8'h3B, 8'h3A, 8'h38, 8'h37, 8'h33, 8'h2E, 8'h2A, 8'h23, 8'h1C, 8'h14, 8'h0B, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h2A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h03, 8'h03, 8'h04, 8'h04, 8'h04, 8'h12, 8'h1D, 8'h27, 8'h30, 8'h39, 8'h3E, 8'h44, 8'h48, 8'h4B, 8'h4D, 8'h4E, 8'h4E, 8'h4D, 8'h4B, 8'h48, 8'h44, 8'h3E, 8'h39, 8'h30, 8'h27, 8'h1D, 8'h12, 8'h04, 8'h04, 8'h04, 8'h03, 8'h03, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2B, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h6C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h62, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h35, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h08, 8'h0B, 8'h0F, 8'h12, 8'h12, 8'h12, 8'h1E, 8'h29, 8'h33, 8'h3B, 8'h43, 8'h49, 8'h4E, 8'h53, 8'h55, 8'h57, 8'h58, 8'h58, 8'h57, 8'h55, 8'h53, 8'h4E, 8'h49, 8'h43, 8'h3B, 8'h33, 8'h29, 8'h1E, 8'h12, 8'h12, 8'h12, 8'h0F, 8'h0B, 8'h08, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h36, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h62, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h11, 8'h1A, 8'h22, 8'h29, 8'h28, 8'h27, 8'h30, 8'h37, 8'h3E, 8'h44, 8'h49, 8'h4D, 8'h51, 8'h54, 8'h56, 8'h58, 8'h58, 8'h58, 8'h58, 8'h56, 8'h54, 8'h51, 8'h4D, 8'h49, 8'h44, 8'h3E, 8'h37, 8'h30, 8'h27, 8'h28, 8'h29, 8'h22, 8'h1A, 8'h11, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h42, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h59, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4F, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0E, 8'h1E, 8'h2C, 8'h39, 8'h44, 8'h43, 8'h41, 8'h44, 8'h48, 8'h4A, 8'h4C, 8'h4E, 8'h50, 8'h51, 8'h53, 8'h53, 8'h54, 8'h54, 8'h54, 8'h54, 8'h53, 8'h53, 8'h51, 8'h50, 8'h4E, 8'h4C, 8'h4A, 8'h48, 8'h44, 8'h41, 8'h43, 8'h44, 8'h39, 8'h2C, 8'h1E, 8'h0E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h4F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h47, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h58, 8'h04, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h02, 8'h03, 8'h04, 8'h04, 8'h16, 8'h29, 8'h3B, 8'h4C, 8'h5A, 8'h58, 8'h55, 8'h54, 8'h54, 8'h53, 8'h52, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h51, 8'h52, 8'h53, 8'h54, 8'h54, 8'h55, 8'h58, 8'h5A, 8'h4C, 8'h3B, 8'h29, 8'h16, 8'h04, 8'h04, 8'h03, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00, 8'h01, 8'h04, 8'h58, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h47, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h40, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5B, 8'h11, 8'h07, 8'h00, 8'h00, 8'h01, 8'h06, 8'h0A, 8'h0F, 8'h12, 8'h11, 8'h22, 8'h35, 8'h46, 8'h56, 8'h63, 8'h62, 8'h5F, 8'h5B, 8'h59, 8'h57, 8'h55, 8'h52, 8'h52, 8'h50, 8'h50, 8'h4F, 8'h4F, 8'h4E, 8'h4E, 8'h4F, 8'h4F, 8'h50, 8'h50, 8'h52, 8'h52, 8'h55, 8'h57, 8'h59, 8'h5B, 8'h5F, 8'h62, 8'h63, 8'h56, 8'h46, 8'h35, 8'h22, 8'h11, 8'h12, 8'h0F, 8'h0A, 8'h06, 8'h01, 8'h00, 8'h00, 8'h07, 8'h11, 8'h5B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h40, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3B, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h58, 8'h27, 8'h0F, 8'h00, 8'h00, 8'h02, 8'h0D, 8'h18, 8'h22, 8'h29, 8'h26, 8'h32, 8'h3F, 8'h4B, 8'h57, 8'h60, 8'h5F, 8'h5D, 8'h59, 8'h58, 8'h55, 8'h54, 8'h51, 8'h50, 8'h4F, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4F, 8'h4F, 8'h50, 8'h51, 8'h54, 8'h55, 8'h58, 8'h59, 8'h5D, 8'h5F, 8'h60, 8'h57, 8'h4B, 8'h3F, 8'h32, 8'h26, 8'h29, 8'h22, 8'h17, 8'h0D, 8'h02, 8'h00, 8'h00, 8'h0F, 8'h27, 8'h58, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h37, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h42, 8'h1A, 8'h00, 8'h00, 8'h04, 8'h16, 8'h28, 8'h39, 8'h44, 8'h41, 8'h45, 8'h4B, 8'h4F, 8'h53, 8'h57, 8'h57, 8'h55, 8'h54, 8'h52, 8'h52, 8'h50, 8'h4F, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h4F, 8'h50, 8'h52, 8'h52, 8'h54, 8'h55, 8'h57, 8'h57, 8'h53, 8'h4F, 8'h4B, 8'h45, 8'h41, 8'h44, 8'h39, 8'h27, 8'h16, 8'h04, 8'h00, 8'h00, 8'h1A, 8'h42, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h37, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h57, 8'h24, 8'h04, 8'h04, 8'h08, 8'h1F, 8'h36, 8'h4C, 8'h5A, 8'h55, 8'h53, 8'h53, 8'h51, 8'h51, 8'h50, 8'h50, 8'h50, 8'h4F, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4F, 8'h50, 8'h50, 8'h50, 8'h51, 8'h51, 8'h53, 8'h53, 8'h55, 8'h5A, 8'h4C, 8'h35, 8'h1F, 8'h08, 8'h04, 8'h04, 8'h24, 8'h57, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h33, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h60, 8'h30, 8'h11, 8'h11, 8'h15, 8'h2B, 8'h41, 8'h56, 8'h63, 8'h5F, 8'h5A, 8'h57, 8'h52, 8'h4F, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4F, 8'h52, 8'h57, 8'h5A, 8'h5F, 8'h63, 8'h56, 8'h40, 8'h2B, 8'h15, 8'h11, 8'h11, 8'h30, 8'h60, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h33, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h5E, 8'h3C, 8'h27, 8'h27, 8'h29, 8'h39, 8'h48, 8'h57, 8'h60, 8'h5D, 8'h58, 8'h55, 8'h51, 8'h4E, 8'h4B, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4B, 8'h4E, 8'h51, 8'h55, 8'h58, 8'h5D, 8'h60, 8'h57, 8'h47, 8'h39, 8'h29, 8'h27, 8'h27, 8'h3C, 8'h5E, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'h37, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h49, 8'h41, 8'h42, 8'h41, 8'h47, 8'h4E, 8'h53, 8'h57, 8'h55, 8'h53, 8'h52, 8'h4F, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4F, 8'h52, 8'h53, 8'h55, 8'h57, 8'h53, 8'h4E, 8'h47, 8'h41, 8'h42, 8'h41, 8'h49, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h37, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h53, 8'h56, 8'h57, 8'h54, 8'h53, 8'h52, 8'h51, 8'h50, 8'h50, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h50, 8'h50, 8'h51, 8'h53, 8'h53, 8'h54, 8'h57, 8'h56, 8'h53, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'h3A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h58, 8'h60, 8'h60, 8'h5D, 8'h58, 8'h54, 8'h4F, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4F, 8'h54, 8'h58, 8'h5D, 8'h60, 8'h60, 8'h58, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3A, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h5D, 8'h5E, 8'h5B, 8'h57, 8'h52, 8'h4E, 8'h4B, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4B, 8'h4E, 8'h53, 8'h57, 8'h5B, 8'h5E, 8'h5D, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h52, 8'h56, 8'h56, 8'h54, 8'h52, 8'h50, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h50, 8'h52, 8'h54, 8'h56, 8'h56, 8'h52, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h50, 8'h50, 8'h4F, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h4F, 8'h50, 8'h50, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hDC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD3, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD0, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC3, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h50, 8'h50, 8'h4F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4F, 8'h50, 8'h50, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4E, 8'h53, 8'h54, 8'h50, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h50, 8'h54, 8'h53, 8'h4E, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4F, 8'h54, 8'h55, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h55, 8'h54, 8'h4F, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h50, 8'h51, 8'h52, 8'h52, 8'h51, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h51, 8'h52, 8'h52, 8'h51, 8'h50, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h53, 8'h4D, 8'h4C, 8'h4F, 8'h57, 8'h50, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h50, 8'h57, 8'h4F, 8'h4C, 8'h4D, 8'h53, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h5E, 8'h56, 8'h45, 8'h44, 8'h4D, 8'h60, 8'h53, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h53, 8'h60, 8'h4D, 8'h44, 8'h45, 8'h56, 8'h5E, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD0, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4E, 8'h60, 8'h55, 8'h3D, 8'h3B, 8'h48, 8'h63, 8'h54, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h54, 8'h63, 8'h48, 8'h3B, 8'h3D, 8'h55, 8'h60, 8'h4E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD3, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h51, 8'h57, 8'h4B, 8'h32, 8'h30, 8'h3D, 8'h59, 8'h53, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h52, 8'h59, 8'h3D, 8'h30, 8'h32, 8'h4B, 8'h57, 8'h51, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h42, 8'h39, 8'h25, 8'h23, 8'h2E, 8'h44, 8'h4E, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h4D, 8'h44, 8'h2E, 8'h23, 8'h25, 8'h39, 8'h42, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5B, 8'h27, 8'h22, 8'h16, 8'h15, 8'h1B, 8'h28, 8'h47, 8'h55, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h55, 8'h47, 8'h28, 8'h1B, 8'h15, 8'h16, 8'h22, 8'h27, 8'h5B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h5C, 8'h11, 8'h0F, 8'h0A, 8'h09, 8'h0C, 8'h12, 8'h40, 8'h57, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h57, 8'h3F, 8'h12, 8'h0C, 8'h09, 8'h0A, 8'h0F, 8'h11, 8'h5C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h52, 8'h04, 8'h03, 8'h02, 8'h02, 8'h03, 8'h04, 8'h35, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h34, 8'h04, 8'h03, 8'h02, 8'h02, 8'h03, 8'h04, 8'h52, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h3E, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h26, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h25, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h17, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h17, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h25, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'h3A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h5B, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h41, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h41, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h5B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3A, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h36, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h36, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'h37, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h37, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h17, 8'h57, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h57, 8'h17, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h39, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h34, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h33, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h2C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0A, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h0A, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2A, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h33, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1E, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h34, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h37, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h16, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h15, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h37, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3B, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h0D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h3B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h40, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h06, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h40, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h40, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h47, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h38, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h39, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h47, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4F, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h33, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h33, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h4F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h59, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h62, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h62, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h26, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h6C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h26, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h26, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h74, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h27, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h7E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h88, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h87, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h92, 8'h43, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h43, 8'h91, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9C, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h9B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA7, 8'h41, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h41, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBE, 8'h3E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3E, 8'hBE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'h3C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'h37, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h37, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'h36, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h35, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h35, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'h33, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h32, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h35, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h33, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h3D, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h3C, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4C, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h4A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5D, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h5C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6E, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h6D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7F, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h7E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8F, 8'h43, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h27, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h43, 8'h8E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9F, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h26, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h27, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h9E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAF, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h27, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h27, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hAE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC0, 8'h3B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h29, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3B, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'h36, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h2D, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h2D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h36, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h31, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h31, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'h2C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h36, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h36, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2C, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'h30, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h55, 8'h05, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3D, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3D, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h05, 8'h55, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h30, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3B, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h45, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h45, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4A, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h13, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h13, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h49, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h59, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h56, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h57, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6C, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h28, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h28, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h46, 8'h6B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h82, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h36, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h15, 8'h57, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h57, 8'h16, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h36, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h80, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h99, 8'h41, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h54, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h54, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h41, 8'h99, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAF, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h03, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h02, 8'h31, 8'h51, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h32, 8'h02, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h03, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'hAF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'h3A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h10, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h09, 8'h3D, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3E, 8'h09, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h10, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3A, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'h34, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h58, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h14, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h14, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h58, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h34, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h2D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h53, 8'h3C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3C, 8'h53, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2D, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h2B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h50, 8'h04, 8'h03, 8'h02, 8'h02, 8'h02, 8'h04, 8'h2E, 8'h56, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h57, 8'h2E, 8'h04, 8'h02, 8'h02, 8'h02, 8'h03, 8'h04, 8'h50, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2B, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'h34, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h5A, 8'h12, 8'h0D, 8'h09, 8'h08, 8'h0B, 8'h11, 8'h39, 8'h59, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h59, 8'h39, 8'h11, 8'h0B, 8'h08, 8'h09, 8'h0D, 8'h12, 8'h5A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h47, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h59, 8'h28, 8'h1F, 8'h13, 8'h12, 8'h18, 8'h27, 8'h43, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h43, 8'h27, 8'h18, 8'h11, 8'h13, 8'h1F, 8'h28, 8'h59, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h46, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h60, 8'h48, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h55, 8'h44, 8'h33, 8'h21, 8'h1F, 8'h29, 8'h42, 8'h4C, 8'h52, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h52, 8'h4C, 8'h42, 8'h29, 8'h1E, 8'h21, 8'h33, 8'h44, 8'h55, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h48, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h79, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h51, 8'h59, 8'h44, 8'h2D, 8'h2A, 8'h37, 8'h57, 8'h53, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h53, 8'h57, 8'h37, 8'h29, 8'h2D, 8'h44, 8'h59, 8'h51, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h77, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h95, 8'h40, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4E, 8'h63, 8'h4F, 8'h38, 8'h36, 8'h42, 8'h60, 8'h56, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h56, 8'h60, 8'h42, 8'h34, 8'h38, 8'h4F, 8'h63, 8'h4E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h40, 8'h93, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h38, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h5F, 8'h51, 8'h41, 8'h40, 8'h48, 8'h5E, 8'h55, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h55, 8'h5E, 8'h48, 8'h3F, 8'h41, 8'h51, 8'h5F, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h38, 8'hB1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h57, 8'h51, 8'h4B, 8'h4A, 8'h4E, 8'h56, 8'h51, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h51, 8'h56, 8'h4E, 8'h49, 8'h4B, 8'h51, 8'h57, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hD0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'h2A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h50, 8'h50, 8'h52, 8'h52, 8'h51, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h51, 8'h52, 8'h52, 8'h50, 8'h50, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2A, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h2E, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4F, 8'h55, 8'h55, 8'h53, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h53, 8'h55, 8'h55, 8'h4F, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h2E, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3A, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4B, 8'h4F, 8'h54, 8'h54, 8'h52, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h52, 8'h54, 8'h54, 8'h4F, 8'h4B, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h39, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4B, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h50, 8'h51, 8'h4F, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4F, 8'h51, 8'h50, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h4A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5E, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h5C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7A, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h79, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9D, 8'h39, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h39, 8'h9C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'h2F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h2F, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'h29, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h29, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h2D, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h2D, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h3A, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h3A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h4B, 8'h49, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h49, 8'h4B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h5F, 8'h46, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h46, 8'h5F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7C, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'h7C, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9E, 8'h35, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h35, 8'h9E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'h29, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h29, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h24, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h24, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'h2E, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h2E, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h48, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h48, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h69, 8'h42, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h42, 8'h69, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h88, 8'h3D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3D, 8'h88, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA6, 8'h38, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h38, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC0, 8'h32, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h32, 8'hC0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'h2D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h2D, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'h30, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h30, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h49, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h49, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h75, 8'h39, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h39, 8'h75, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h2B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h2B, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h24, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h24, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h2C, 8'h4B, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4B, 8'h2C, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'h44, 8'h45, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h45, 8'h43, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h63, 8'h3F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h3F, 8'h62, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h81, 8'h39, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h39, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9F, 8'h36, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h36, 8'h9D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h35, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h34, 8'hB9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h34, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h34, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'h3B, 8'h47, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h47, 8'h3B, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h55, 8'h3F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3F, 8'h54, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h80, 8'h33, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h33, 8'h7F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB3, 8'h24, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h24, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h21, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h21, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h38, 8'h43, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h43, 8'h38, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h68, 8'h35, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h35, 8'h68, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA6, 8'h22, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h22, 8'hA6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'h1B, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h1B, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h2D, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h2D, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h57, 8'h38, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h38, 8'h57, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h8D, 8'h27, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h27, 8'h8D, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBB, 8'h1F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h1F, 8'hBB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h2C, 8'h47, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h47, 8'h2C, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'h4F, 8'h3A, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3A, 8'h4F, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'h7B, 8'h29, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h51, 8'h29, 8'h7B, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hA3, 8'h22, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h22, 8'hA3, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC1, 8'h2E, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h48, 8'h2E, 8'hC1, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h4E, 8'h39, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h3A, 8'h4E, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h76, 8'h28, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h29, 8'h76, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'h9B, 8'h21, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h21, 8'h9B, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hB9, 8'h2E, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h2F, 8'hB9, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'h50, 8'h36, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h36, 8'h50, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE2, 8'h7C, 8'h24, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h24, 8'h7C, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hA2, 8'h1C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h1C, 8'hA2, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC1, 8'h2D, 8'h44, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h44, 8'h2D, 8'hC1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'h57, 8'h33, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h33, 8'h57, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'h8D, 8'h1F, 8'h4C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4C, 8'h1F, 8'h8D, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBB, 8'h17, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h17, 8'hBB, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hDA, 8'h2D, 8'h41, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h41, 8'h2D, 8'hDA, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'h5F, 8'h32, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h32, 8'h5F, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hA0, 8'h21, 8'h46, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h46, 8'h21, 8'hA0, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hD5, 8'h1B, 8'h43, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h43, 8'h1B, 8'hD5, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF6, 8'h32, 8'h3F, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h3F, 8'h32, 8'hF6, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h63, 8'h3B, 8'h40, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h40, 8'h3B, 8'h63, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA3, 8'h37, 8'h36, 8'h50, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h50, 8'h36, 8'h38, 8'hA3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'h3B, 8'h31, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h31, 8'h3C, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'h53, 8'h38, 8'h44, 8'h4C, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4C, 8'h44, 8'h39, 8'h54, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h7E, 8'h4C, 8'h34, 8'h4C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4C, 8'h34, 8'h4D, 8'h7E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB2, 8'h67, 8'h20, 8'h4A, 8'h4F, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4F, 8'h4A, 8'h1F, 8'h67, 8'hB3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'h80, 8'h19, 8'h48, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h48, 8'h18, 8'h81, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h9C, 8'h2F, 8'h41, 8'h49, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h49, 8'h41, 8'h2E, 8'h9D, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB7, 8'h61, 8'h37, 8'h40, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h40, 8'h37, 8'h60, 8'hB8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hA1, 8'h2B, 8'h36, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h36, 8'h2B, 8'hA1, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'hD6, 8'h29, 8'h31, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h31, 8'h29, 8'hD6, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'h40, 8'h3A, 8'h44, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h44, 8'h3A, 8'h40, 8'hF6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h6F, 8'h50, 8'h33, 8'h46, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h46, 8'h33, 8'h50, 8'h6F, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA9, 8'h6D, 8'h1E, 8'h3F, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h3F, 8'h1E, 8'h6D, 8'hA9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'h88, 8'h16, 8'h3C, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h3C, 8'h16, 8'h88, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hA4, 8'h2D, 8'h3E, 8'h44, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h44, 8'h3E, 8'h2D, 8'hA4, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBE, 8'h5F, 8'h46, 8'h34, 8'h46, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h46, 8'h33, 8'h46, 8'h5F, 8'hBE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'hA0, 8'h50, 8'h1F, 8'h41, 8'h50, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h50, 8'h41, 8'h1F, 8'h50, 8'hA0, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hD5, 8'h5F, 8'h18, 8'h3E, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h3E, 8'h17, 8'h5F, 8'hD5, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'h79, 8'h2E, 8'h3F, 8'h44, 8'h4A, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4A, 8'h44, 8'h3F, 8'h2D, 8'h79, 8'hF6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h9B, 8'h60, 8'h45, 8'h33, 8'h43, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h43, 8'h33, 8'h45, 8'h60, 8'h9B, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'hA1, 8'h4D, 8'h1E, 8'h3C, 8'h4F, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h4F, 8'h3C, 8'h1E, 8'h4D, 8'hA0, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hD6, 8'h5A, 8'h16, 8'h38, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h38, 8'h16, 8'h5A, 8'hD5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF6, 8'h73, 8'h2D, 8'h3E, 8'h43, 8'h48, 8'h4B, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4B, 8'h48, 8'h43, 8'h3E, 8'h2D, 8'h73, 8'hF6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h97, 8'h5F, 8'h4C, 8'h33, 8'h3D, 8'h48, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h48, 8'h3D, 8'h33, 8'h4D, 8'h5F, 8'h97, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC1, 8'hA0, 8'h60, 8'h1F, 8'h30, 8'h43, 8'h50, 8'h4F, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4F, 8'h50, 8'h43, 8'h30, 8'h1F, 8'h61, 8'hA0, 8'hC1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE4, 8'hD5, 8'h74, 8'h18, 8'h2B, 8'h40, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h40, 8'h2B, 8'h18, 8'h76, 8'hD5, 8'hE4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF6, 8'h8F, 8'h2E, 8'h3B, 8'h3F, 8'h44, 8'h48, 8'h4A, 8'h4D, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4D, 8'h4A, 8'h48, 8'h44, 8'h3F, 8'h3B, 8'h2E, 8'h90, 8'hF6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h60, 8'h5C, 8'h41, 8'h33, 8'h3D, 8'h45, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4F, 8'h4D, 8'h45, 8'h3D, 8'h33, 8'h41, 8'h5C, 8'h60, 8'hAE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hA1, 8'h87, 8'h43, 8'h1E, 8'h30, 8'h40, 8'h4D, 8'h50, 8'h4F, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4F, 8'h50, 8'h4D, 8'h40, 8'h30, 8'h1E, 8'h43, 8'h87, 8'hA1, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hD6, 8'hAC, 8'h4C, 8'h16, 8'h2B, 8'h3C, 8'h4B, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4B, 8'h3C, 8'h2B, 8'h16, 8'h4C, 8'hAC, 8'hD6, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF6, 8'hC9, 8'h65, 8'h2D, 8'h3A, 8'h3F, 8'h42, 8'h45, 8'h48, 8'h4A, 8'h4C, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4B, 8'h4A, 8'h48, 8'h46, 8'h42, 8'h3F, 8'h3B, 8'h2D, 8'h65, 8'hC9, 8'hF6, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'h8B, 8'h5F, 8'h5B, 8'h47, 8'h34, 8'h36, 8'h3D, 8'h43, 8'h48, 8'h4C, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h4F, 8'h4C, 8'h48, 8'h43, 8'h3D, 8'h36, 8'h34, 8'h48, 8'h5C, 8'h5F, 8'h8B, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hBA, 8'hA0, 8'h86, 8'h52, 8'h23, 8'h24, 8'h30, 8'h3B, 8'h45, 8'h4C, 8'h50, 8'h50, 8'h50, 8'h50, 8'h4F, 8'h4F, 8'h4F, 8'h4F, 8'h50, 8'h50, 8'h50, 8'h50, 8'h4C, 8'h43, 8'h3B, 8'h30, 8'h23, 8'h23, 8'h53, 8'h87, 8'hA0, 8'hBA, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hE1, 8'hD5, 8'hAB, 8'h61, 8'h1E, 8'h1E, 8'h2B, 8'h37, 8'h42, 8'h49, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4D, 8'h4D, 8'h4D, 8'h4D, 8'h4E, 8'h4E, 8'h4E, 8'h4E, 8'h49, 8'h40, 8'h37, 8'h2B, 8'h1C, 8'h1E, 8'h62, 8'hAC, 8'hD5, 8'hE1, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF8, 8'hF6, 8'hC8, 8'h7A, 8'h35, 8'h34, 8'h3A, 8'h3E, 8'h41, 8'h42, 8'h44, 8'h45, 8'h46, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h46, 8'h45, 8'h44, 8'h42, 8'h40, 8'h3E, 8'h3B, 8'h32, 8'h35, 8'h7C, 8'hC9, 8'hF6, 8'hF8, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h9C, 8'h65, 8'h65, 8'h5B, 8'h4E, 8'h42, 8'h37, 8'h33, 8'h35, 8'h38, 8'h3A, 8'h3B, 8'h3B, 8'h3B, 8'h3B, 8'h3A, 8'h38, 8'h35, 8'h33, 8'h37, 8'h42, 8'h4F, 8'h5C, 8'h63, 8'h65, 8'h9E, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hC5, 8'hA4, 8'hA3, 8'h86, 8'h63, 8'h45, 8'h2A, 8'h1E, 8'h23, 8'h28, 8'h2B, 8'h2C, 8'h2D, 8'h2D, 8'h2C, 8'h2B, 8'h28, 8'h23, 8'h1F, 8'h2A, 8'h45, 8'h64, 8'h87, 8'hA3, 8'hA4, 8'hC5, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hE5, 8'hD7, 8'hD7, 8'hAB, 8'h79, 8'h4D, 8'h27, 8'h16, 8'h1C, 8'h22, 8'h26, 8'h27, 8'h28, 8'h28, 8'h27, 8'h26, 8'h22, 8'h1C, 8'h17, 8'h27, 8'h4E, 8'h7A, 8'hAC, 8'hD6, 8'hD7, 8'hE6, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF9, 8'hF6, 8'hF6, 8'hC8, 8'h93, 8'h66, 8'h3E, 8'h2D, 8'h32, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h39, 8'h32, 8'h2D, 8'h3E, 8'h67, 8'h95, 8'hC9, 8'hF6, 8'hF6, 8'hF9, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hB1, 8'h8C, 8'h6D, 8'h5F, 8'h63, 8'h68, 8'h64, 8'h60, 8'h5F, 8'h5F, 8'h60, 8'h64, 8'h68, 8'h63, 8'h5F, 8'h6D, 8'h8D, 8'hB2, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hD0, 8'hBB, 8'hA8, 8'hA0, 8'hA3, 8'hA6, 8'h9A, 8'h93, 8'h8F, 8'h8F, 8'h93, 8'h9A, 8'hA6, 8'hA3, 8'hA0, 8'hA8, 8'hBC, 8'hD1, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hEB, 8'hE1, 8'hD9, 8'hD5, 8'hD6, 8'hD8, 8'hC8, 8'hBD, 8'hB8, 8'hB8, 8'hBD, 8'hC8, 8'hD8, 8'hD6, 8'hD5, 8'hD9, 8'hE1, 8'hEB, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFA, 8'hF8, 8'hF7, 8'hF6, 8'hF6, 8'hF6, 8'hE6, 8'hDB, 8'hD6, 8'hD6, 8'hDB, 8'hE6, 8'hF6, 8'hF6, 8'hF6, 8'hF7, 8'hF8, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hE9, 8'hE5, 8'hE5, 8'hE9, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hF2, 8'hF0, 8'hF0, 8'hF2, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF9, 8'hF8, 8'hF8, 8'hF9, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF}; 
reg	[7:0]	pattern_data_G1 [0:39999] = '{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFD, 8'hFD, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hFB, 8'hFB, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF9, 8'hF7, 8'hF7, 8'hF9, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFD, 8'hFD, 8'hFC, 8'hFC, 8'hFD, 8'hF8, 8'hF5, 8'hF3, 8'hF3, 8'hF5, 8'hF8, 8'hFD, 8'hFC, 8'hFC, 8'hFD, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF9, 8'hF6, 8'hF4, 8'hF3, 8'hF3, 8'hF4, 8'hEF, 8'hEC, 8'hEA, 8'hEA, 8'hEC, 8'hEF, 8'hF4, 8'hF3, 8'hF3, 8'hF4, 8'hF6, 8'hF9, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hF2, 8'hEB, 8'hE6, 8'hE3, 8'hE4, 8'hE5, 8'hE2, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hE2, 8'hE5, 8'hE4, 8'hE3, 8'hE6, 8'hEB, 8'hF2, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE8, 8'hDE, 8'hD5, 8'hD0, 8'hD2, 8'hD4, 8'hD2, 8'hD1, 8'hD0, 8'hD0, 8'hD1, 8'hD2, 8'hD4, 8'hD2, 8'hD0, 8'hD5, 8'hDE, 8'hE8, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFC, 8'hFC, 8'hEE, 8'hE0, 8'hD3, 8'hC8, 8'hC1, 8'hC4, 8'hC6, 8'hC6, 8'hC5, 8'hC6, 8'hC6, 8'hC5, 8'hC6, 8'hC6, 8'hC4, 8'hC1, 8'hC8, 8'hD3, 8'hE0, 8'hEE, 8'hFC, 8'hFC, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF7, 8'hF3, 8'hF3, 8'hE6, 8'hD8, 8'hCB, 8'hC1, 8'hBB, 8'hBD, 8'hC0, 8'hC0, 8'hC0, 8'hC1, 8'hC1, 8'hC0, 8'hC0, 8'hC0, 8'hBD, 8'hBB, 8'hC1, 8'hCB, 8'hD8, 8'hE6, 8'hF3, 8'hF4, 8'hF7, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hEE, 8'hE5, 8'hE5, 8'hDC, 8'hD2, 8'hC9, 8'hC2, 8'hBD, 8'hBF, 8'hC1, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC1, 8'hBF, 8'hBD, 8'hC2, 8'hC9, 8'hD2, 8'hDC, 8'hE4, 8'hE5, 8'hEE, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE2, 8'hD2, 8'hD2, 8'hCF, 8'hCC, 8'hC8, 8'hC5, 8'hC4, 8'hC5, 8'hC6, 8'hC6, 8'hC6, 8'hC7, 8'hC7, 8'hC6, 8'hC6, 8'hC6, 8'hC5, 8'hC4, 8'hC5, 8'hC8, 8'hCC, 8'hCF, 8'hD2, 8'hD3, 8'hE2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFC, 8'hEE, 8'hD8, 8'hC4, 8'hC4, 8'hC6, 8'hC7, 8'hC8, 8'hC9, 8'hC9, 8'hC9, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hC9, 8'hC9, 8'hC9, 8'hC8, 8'hC7, 8'hC6, 8'hC4, 8'hC5, 8'hD8, 8'hEF, 8'hFC, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF6, 8'hF3, 8'hE6, 8'hD1, 8'hBE, 8'hBE, 8'hC2, 8'hC5, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC5, 8'hC2, 8'hBD, 8'hBE, 8'hD1, 8'hE7, 8'hF3, 8'hF6, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hEB, 8'hE3, 8'hDC, 8'hCD, 8'hBF, 8'hC0, 8'hC4, 8'hC6, 8'hC9, 8'hCB, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCB, 8'hC9, 8'hC6, 8'hC4, 8'hBF, 8'hC0, 8'hCD, 8'hDC, 8'hE3, 8'hEB, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDE, 8'hD1, 8'hCF, 8'hCA, 8'hC4, 8'hC5, 8'hC7, 8'hC9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC9, 8'hC7, 8'hC5, 8'hC4, 8'hCA, 8'hD0, 8'hD1, 8'hDE, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hEF, 8'hD3, 8'hC2, 8'hC6, 8'hC8, 8'hC8, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hC9, 8'hC8, 8'hC8, 8'hC6, 8'hC2, 8'hD3, 8'hF0, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF3, 8'hE7, 8'hCB, 8'hBB, 8'hC2, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hC2, 8'hBB, 8'hCB, 8'hE7, 8'hF3, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hE4, 8'hDC, 8'hC9, 8'hBE, 8'hC4, 8'hC8, 8'hCB, 8'hCD, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCD, 8'hCB, 8'hC8, 8'hC4, 8'hBE, 8'hC9, 8'hDC, 8'hE4, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hD1, 8'hD0, 8'hC8, 8'hC3, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hC3, 8'hC8, 8'hCF, 8'hD1, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hDE, 8'hC3, 8'hC6, 8'hC8, 8'hC8, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hC8, 8'hC8, 8'hC5, 8'hC3, 8'hDE, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hF3, 8'hD7, 8'hBC, 8'hC2, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC1, 8'hBC, 8'hD7, 8'hF3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hE4, 8'hD1, 8'hBE, 8'hC4, 8'hC9, 8'hCC, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCC, 8'hC9, 8'hC2, 8'hBE, 8'hD1, 8'hE4, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'hD1, 8'hCB, 8'hC4, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hC4, 8'hCB, 8'hD1, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hD6, 8'hC3, 8'hC7, 8'hC8, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hC8, 8'hC7, 8'hC3, 8'hD6, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hF3, 8'hCE, 8'hBC, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC5, 8'hBC, 8'hCE, 8'hF3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hE4, 8'hCB, 8'hBE, 8'hC6, 8'hCC, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCC, 8'hC6, 8'hBE, 8'hCB, 8'hE4, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE1, 8'hD1, 8'hC9, 8'hC4, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC4, 8'hC9, 8'hD1, 8'hE1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hD7, 8'hC3, 8'hC8, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC8, 8'hC3, 8'hD7, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF3, 8'hD0, 8'hBC, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hBC, 8'hD0, 8'hF3, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE3, 8'hCC, 8'hBE, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hBE, 8'hCC, 8'hE3, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'hD1, 8'hC8, 8'hC4, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC4, 8'hC8, 8'hD1, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE5, 8'hC2, 8'hC6, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC6, 8'hC2, 8'hE5, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDD, 8'hBB, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hBB, 8'hDD, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'hD5, 8'hBE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hBE, 8'hD5, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hCC, 8'hC3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC3, 8'hCC, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hC8, 8'hC6, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC6, 8'hC8, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF3, 8'hC1, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hC1, 8'hF3, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hE3, 8'hC2, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hC2, 8'hE3, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hD1, 8'hC5, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC5, 8'hD1, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE2, 8'hC2, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hC2, 8'hE2, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hDA, 8'hBB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBB, 8'hDA, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hD2, 8'hBE, 8'hCB, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCB, 8'hBE, 8'hD2, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hCB, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hCB, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hCE, 8'hC5, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC5, 8'hCE, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC7, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hC7, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC5, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hC5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC7, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC7, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC4, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hC4, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF3, 8'hBE, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCD, 8'hCD, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hBE, 8'hF3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE3, 8'hBF, 8'hC9, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCE, 8'hCF, 8'hCF, 8'hCE, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC9, 8'hBF, 8'hE3, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD1, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCA, 8'hCA, 8'hC9, 8'hC9, 8'hCD, 8'hCF, 8'hD1, 8'hD1, 8'hCF, 8'hCD, 8'hC9, 8'hC9, 8'hCA, 8'hCA, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hD1, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF4, 8'hC2, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCF, 8'hD1, 8'hD3, 8'hD3, 8'hD1, 8'hCF, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC2, 8'hF4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hEA, 8'hBB, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCD, 8'hCF, 8'hD1, 8'hD1, 8'hD1, 8'hD3, 8'hD4, 8'hD4, 8'hD4, 8'hD4, 8'hD3, 8'hD1, 8'hD1, 8'hD1, 8'hCF, 8'hCD, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hBB, 8'hEA, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hDD, 8'hBE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hD1, 8'hD6, 8'hDB, 8'hDC, 8'hDC, 8'hDA, 8'hD6, 8'hD5, 8'hD5, 8'hD6, 8'hDA, 8'hDC, 8'hDC, 8'hDA, 8'hD6, 8'hD1, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBE, 8'hDD, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hCE, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hC9, 8'hCB, 8'hD5, 8'hDF, 8'hE7, 8'hEB, 8'hEB, 8'hE1, 8'hD9, 8'hD4, 8'hD4, 8'hD9, 8'hE1, 8'hEB, 8'hEB, 8'hE7, 8'hDF, 8'hD5, 8'hCB, 8'hC9, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hCE, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hED, 8'hC2, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCA, 8'hCD, 8'hD8, 8'hE2, 8'hEB, 8'hEE, 8'hED, 8'hE0, 8'hD4, 8'hCD, 8'hCD, 8'hD4, 8'hE0, 8'hED, 8'hEE, 8'hEA, 8'hE2, 8'hD8, 8'hCD, 8'hCA, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC2, 8'hED, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE4, 8'hBD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCE, 8'hD0, 8'hD3, 8'hD6, 8'hD9, 8'hDB, 8'hD9, 8'hD4, 8'hC7, 8'hBB, 8'hB4, 8'hB4, 8'hBB, 8'hC7, 8'hD4, 8'hD9, 8'hDA, 8'hD9, 8'hD6, 8'hD4, 8'hD0, 8'hCE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBD, 8'hE4, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hD9, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD3, 8'hDB, 8'hDE, 8'hCF, 8'hC3, 8'hB8, 8'hAC, 8'hA2, 8'h99, 8'h91, 8'h8C, 8'h8C, 8'h91, 8'h99, 8'hA2, 8'hAC, 8'hB8, 8'hC3, 8'hCF, 8'hDE, 8'hDB, 8'hD3, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hD9, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hCD, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hCB, 8'hD9, 8'hE8, 8'hEA, 8'hC6, 8'hA6, 8'h8B, 8'h73, 8'h63, 8'h60, 8'h5D, 8'h5B, 8'h5B, 8'h5D, 8'h60, 8'h63, 8'h73, 8'h8B, 8'hA7, 8'hC6, 8'hEC, 8'hE8, 8'hD9, 8'hCB, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hCC, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hEA, 8'hC3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCD, 8'hDC, 8'hEC, 8'hEC, 8'hB9, 8'h8C, 8'h66, 8'h46, 8'h31, 8'h33, 8'h34, 8'h35, 8'h35, 8'h34, 8'h33, 8'h31, 8'h46, 8'h67, 8'h8D, 8'hB9, 8'hEE, 8'hEC, 8'hDC, 8'hCD, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC3, 8'hEA, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hE1, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hD0, 8'hD3, 8'hD6, 8'hDB, 8'hD3, 8'hA0, 8'h73, 8'h4D, 8'h2E, 8'h1A, 8'h1E, 8'h21, 8'h23, 8'h23, 8'h21, 8'h1E, 8'h1A, 8'h2E, 8'h4E, 8'h74, 8'hA0, 8'hD5, 8'hDB, 8'hD6, 8'hD3, 8'hD0, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hE1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD7, 8'hC1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hD9, 8'hDE, 8'hC9, 8'hB7, 8'hA2, 8'h7E, 8'h5E, 8'h43, 8'h2D, 8'h1E, 8'h23, 8'h25, 8'h27, 8'h27, 8'h25, 8'h23, 8'h1E, 8'h2D, 8'h43, 8'h5E, 8'h7E, 8'hA3, 8'hB7, 8'hC9, 8'hDE, 8'hD9, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC1, 8'hD7, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hCC, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hCF, 8'hE3, 8'hEA, 8'hB7, 8'h88, 8'h63, 8'h55, 8'h49, 8'h3D, 8'h35, 8'h2F, 8'h32, 8'h34, 8'h34, 8'h34, 8'h34, 8'h32, 8'h2F, 8'h35, 8'h3E, 8'h49, 8'h55, 8'h63, 8'h89, 8'hB8, 8'hEA, 8'hE3, 8'hCF, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hCC, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hD1, 8'hE7, 8'hEC, 8'hA5, 8'h61, 8'h32, 8'h36, 8'h39, 8'h3A, 8'h3D, 8'h3C, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3C, 8'h3D, 8'h3A, 8'h38, 8'h36, 8'h32, 8'h62, 8'hA5, 8'hEC, 8'hE7, 8'hD1, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC3, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE4, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hD4, 8'hDA, 8'hD3, 8'h8C, 8'h48, 8'h1B, 8'h27, 8'h32, 8'h39, 8'h41, 8'h44, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h44, 8'h41, 8'h39, 8'h31, 8'h27, 8'h1A, 8'h49, 8'h8D, 8'hD3, 8'hDA, 8'hD4, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hE4, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hD9, 8'hC1, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hDB, 8'hD8, 8'hBE, 8'hA2, 8'h6F, 8'h3F, 8'h1F, 8'h2B, 8'h35, 8'h3C, 8'h43, 8'h46, 8'h48, 8'h47, 8'h47, 8'h47, 8'h47, 8'h48, 8'h46, 8'h43, 8'h3C, 8'h34, 8'h2B, 8'h1F, 8'h40, 8'h70, 8'hA2, 8'hBE, 8'hD9, 8'hDB, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC1, 8'hD9, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hCC, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCE, 8'hE7, 8'hDD, 8'h99, 8'h64, 8'h4F, 8'h3B, 8'h30, 8'h37, 8'h3C, 8'h40, 8'h44, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h44, 8'h40, 8'h3C, 8'h37, 8'h2F, 8'h3C, 8'h4F, 8'h64, 8'h99, 8'hDE, 8'hE7, 8'hCE, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hCC, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hEC, 8'hD9, 8'h7A, 8'h33, 8'h36, 8'h3A, 8'h3D, 8'h40, 8'h42, 8'h43, 8'h45, 8'h45, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h45, 8'h45, 8'h43, 8'h42, 8'h40, 8'h3C, 8'h3A, 8'h36, 8'h33, 8'h7A, 8'hDB, 8'hEC, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hBE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hD4, 8'hDD, 8'hBF, 8'h60, 8'h1C, 8'h2B, 8'h3A, 8'h44, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h44, 8'h3A, 8'h2B, 8'h1C, 8'h60, 8'hC1, 8'hDD, 8'hD4, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBE, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'hC0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD7, 8'hDA, 8'hBD, 8'h92, 8'h50, 8'h20, 8'h2F, 8'h3D, 8'h46, 8'h47, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h47, 8'h46, 8'h3D, 8'h2F, 8'h20, 8'h50, 8'h94, 8'hBD, 8'hDB, 8'hD7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC0, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hE1, 8'hE2, 8'h92, 8'h5B, 8'h43, 8'h30, 8'h38, 8'h40, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h40, 8'h38, 8'h30, 8'h43, 8'h5B, 8'h92, 8'hE2, 8'hE1, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hE5, 8'hE0, 8'h6F, 8'h2F, 8'h39, 8'h3D, 8'h41, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h41, 8'h3D, 8'h39, 8'h2F, 8'h6F, 8'hE1, 8'hE5, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC2, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'hDB, 8'hC7, 8'h55, 8'h1B, 8'h35, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h35, 8'h1B, 8'h55, 8'hC7, 8'hDB, 8'hD1, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBD, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCE, 8'hDC, 8'hC5, 8'h98, 8'h48, 8'h20, 8'h38, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h38, 8'h20, 8'h48, 8'h99, 8'hC5, 8'hDC, 8'hCE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD0, 8'hEB, 8'hA8, 8'h5E, 8'h40, 8'h31, 8'h3D, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h3D, 8'h31, 8'h40, 8'h5E, 8'hA8, 8'hEB, 8'hD1, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC6, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD2, 8'hEE, 8'h8D, 8'h31, 8'h39, 8'h3E, 8'h42, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h42, 8'h3E, 8'h39, 8'h31, 8'h8D, 8'hEE, 8'hD3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCE, 8'hD5, 8'hD9, 8'h74, 8'h1C, 8'h37, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h37, 8'h1C, 8'h74, 8'hD9, 8'hD6, 8'hCE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hC0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD4, 8'hD9, 8'hAC, 8'h5D, 8'h20, 8'h3A, 8'h47, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h47, 8'h3A, 8'h20, 8'h5D, 8'hAD, 8'hD9, 8'hD4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC0, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDC, 8'hDC, 8'h74, 8'h46, 8'h31, 8'h3F, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3F, 8'h31, 8'h46, 8'h74, 8'hDC, 8'hDC, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hCE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hE0, 8'hD8, 8'h46, 8'h35, 8'h3E, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h3E, 8'h35, 8'h47, 8'hD7, 8'hE0, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hCE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD0, 8'hDB, 8'hBE, 8'h2E, 8'h2E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h2E, 8'h2F, 8'hBD, 8'hDB, 8'hD0, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hDA, 8'hCE, 8'h91, 8'h2C, 8'h32, 8'h47, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h47, 8'h32, 8'h2C, 8'h91, 8'hCE, 8'hDA, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC5, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE6, 8'hBD, 8'h5A, 8'h33, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3A, 8'h34, 8'h59, 8'hBD, 8'hE6, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hEB, 8'hAA, 8'h2F, 8'h3A, 8'h41, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h41, 8'h3A, 8'h2F, 8'hAA, 8'hEB, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD0, 8'hE0, 8'h8F, 8'h1B, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3E, 8'h1B, 8'h8F, 8'hE0, 8'hD0, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hDC, 8'hC6, 8'h6E, 8'h20, 8'h41, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h41, 8'h20, 8'h6E, 8'hC6, 8'hDC, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hEA, 8'hA4, 8'h4A, 8'h31, 8'h43, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h43, 8'h31, 8'h4A, 8'hA4, 8'hEA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC2, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hF0, 8'h85, 8'h2D, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3E, 8'h2D, 8'h85, 8'hF0, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC2, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD0, 8'hE2, 8'h6A, 8'h22, 8'h45, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h45, 8'h22, 8'h6A, 8'hE2, 8'hD0, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hDB, 8'hC2, 8'h54, 8'h28, 8'h47, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h47, 8'h28, 8'h54, 8'hC2, 8'hDB, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hEA, 8'h98, 8'h40, 8'h35, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h35, 8'h40, 8'h98, 8'hEA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hCA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hEF, 8'h74, 8'h30, 8'h40, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h40, 8'h30, 8'h74, 8'hEF, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hCA, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hE2, 8'h59, 8'h2B, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2B, 8'h59, 8'hE2, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDA, 8'hC2, 8'h48, 8'h30, 8'h48, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h48, 8'h30, 8'h48, 8'hC2, 8'hDA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE6, 8'h9A, 8'h3B, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3A, 8'h3B, 8'h9A, 8'hE6, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hEC, 8'h76, 8'h32, 8'h42, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h42, 8'h32, 8'h76, 8'hEC, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hE3, 8'h5A, 8'h2F, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2F, 8'h5A, 8'hE3, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD5, 8'hCC, 8'h48, 8'h34, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h34, 8'h48, 8'hCC, 8'hD5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDD, 8'hAC, 8'h3A, 8'h3C, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3C, 8'h3A, 8'hAC, 8'hDD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE3, 8'h8F, 8'h2F, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h2F, 8'h8F, 8'hE3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hE0, 8'h73, 8'h2C, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2C, 8'h73, 8'hE0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hD7, 8'h59, 8'h31, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h47, 8'h47, 8'h46, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h47, 8'h47, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h31, 8'h59, 8'hD7, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD2, 8'hC9, 8'h3F, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h47, 8'h48, 8'h48, 8'h48, 8'h48, 8'h46, 8'h45, 8'h45, 8'h47, 8'h48, 8'h48, 8'h48, 8'h48, 8'h47, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3A, 8'h3F, 8'hC9, 8'hD2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD5, 8'hB9, 8'h2B, 8'h41, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h47, 8'h47, 8'h46, 8'h44, 8'h43, 8'h43, 8'h45, 8'h46, 8'h47, 8'h47, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h41, 8'h2B, 8'hB9, 8'hD5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD9, 8'h9E, 8'h24, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h44, 8'h41, 8'h3F, 8'h3E, 8'h3E, 8'h3E, 8'h3D, 8'h3B, 8'h3B, 8'h3B, 8'h3C, 8'h3D, 8'h3E, 8'h3E, 8'h3E, 8'h40, 8'h41, 8'h44, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h24, 8'h9E, 8'hD9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDD, 8'h7B, 8'h2A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h41, 8'h3A, 8'h35, 8'h31, 8'h2E, 8'h2E, 8'h2E, 8'h2D, 8'h2D, 8'h2D, 8'h2D, 8'h2E, 8'h2E, 8'h2E, 8'h31, 8'h35, 8'h3A, 8'h41, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2A, 8'h7B, 8'hDD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hE2, 8'h52, 8'h37, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h48, 8'h48, 8'h3D, 8'h31, 8'h27, 8'h20, 8'h1C, 8'h1C, 8'h1B, 8'h1A, 8'h1D, 8'h1D, 8'h1B, 8'h1B, 8'h1C, 8'h1C, 8'h20, 8'h28, 8'h31, 8'h3D, 8'h48, 8'h48, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h37, 8'h52, 8'hE2, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE0, 8'h32, 8'h40, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h3A, 8'h2D, 8'h23, 8'h1B, 8'h15, 8'h15, 8'h15, 8'h15, 8'h18, 8'h18, 8'h15, 8'h15, 8'h15, 8'h15, 8'h1B, 8'h23, 8'h2D, 8'h3A, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h40, 8'h32, 8'hE0, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hCE, 8'h23, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h45, 8'h41, 8'h3E, 8'h3D, 8'h39, 8'h34, 8'h32, 8'h30, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h30, 8'h30, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h30, 8'h32, 8'h34, 8'h38, 8'h3D, 8'h3E, 8'h41, 8'h45, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h23, 8'hCE, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD7, 8'hAC, 8'h26, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h45, 8'h3A, 8'h31, 8'h2E, 8'h38, 8'h46, 8'h53, 8'h5E, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h62, 8'h62, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5E, 8'h53, 8'h46, 8'h38, 8'h2E, 8'h31, 8'h3A, 8'h45, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h26, 8'hAC, 8'hD7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'h83, 8'h30, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h48, 8'h44, 8'h32, 8'h20, 8'h1B, 8'h38, 8'h5E, 8'h7E, 8'h99, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA2, 8'hA2, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'h99, 8'h7E, 8'h5E, 8'h37, 8'h1B, 8'h20, 8'h32, 8'h45, 8'h48, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h30, 8'h83, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE6, 8'h60, 8'h39, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h42, 8'h2E, 8'h1B, 8'h15, 8'h3F, 8'h75, 8'hA4, 8'hCA, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD6, 8'hD6, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hCA, 8'hA3, 8'h75, 8'h3E, 8'h15, 8'h1B, 8'h2E, 8'h43, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h39, 8'h60, 8'hE6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE3, 8'h47, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h43, 8'h3E, 8'h3A, 8'h35, 8'h30, 8'h2C, 8'h59, 8'h91, 8'hC2, 8'hE9, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hE9, 8'hC1, 8'h91, 8'h58, 8'h2C, 8'h2F, 8'h35, 8'h3B, 8'h3E, 8'h43, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h47, 8'hE3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h3B, 8'h42, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h40, 8'h31, 8'h2D, 8'h46, 8'h5D, 8'h5F, 8'h82, 8'hAF, 8'hD6, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hD5, 8'hAF, 8'h81, 8'h5F, 8'h5C, 8'h46, 8'h2D, 8'h31, 8'h40, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h42, 8'h3B, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC8, 8'h33, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h49, 8'h3B, 8'h20, 8'h1D, 8'h5D, 8'h97, 8'hA0, 8'hB5, 8'hD0, 8'hE6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hE6, 8'hD0, 8'hB5, 8'hA0, 8'h96, 8'h5D, 8'h1D, 8'h20, 8'h3B, 8'h49, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h33, 8'hC7, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hB7, 8'h2E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h38, 8'h1B, 8'h19, 8'h75, 8'hC7, 8'hD5, 8'hDE, 8'hEA, 8'hF4, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF4, 8'hEA, 8'hDE, 8'hD5, 8'hC7, 8'h75, 8'h18, 8'h1B, 8'h38, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h2E, 8'hB6, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h9F, 8'h2E, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h43, 8'h3F, 8'h38, 8'h2F, 8'h31, 8'h91, 8'hE7, 8'hF6, 8'hF8, 8'hFA, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFA, 8'hF8, 8'hF6, 8'hE6, 8'h91, 8'h30, 8'h2E, 8'h37, 8'h3F, 8'h43, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2E, 8'h9D, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDB, 8'h82, 8'h32, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h40, 8'h2F, 8'h3A, 8'h5A, 8'h63, 8'hAF, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hAF, 8'h62, 8'h5A, 8'h39, 8'h2F, 8'h40, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h32, 8'h80, 8'hDB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE2, 8'h60, 8'h3A, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h48, 8'h3C, 8'h1C, 8'h3D, 8'h93, 8'hA2, 8'hCF, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hCF, 8'hA2, 8'h92, 8'h3C, 8'h1C, 8'h3C, 8'h48, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3A, 8'h60, 8'hE3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE6, 8'h45, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h39, 8'h15, 8'h47, 8'hC2, 8'hD6, 8'hEA, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hEA, 8'hD6, 8'hC1, 8'h45, 8'h15, 8'h39, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h45, 8'hE7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'h35, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h37, 8'h2C, 8'h60, 8'hE1, 8'hF6, 8'hFA, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFA, 8'hF6, 8'hE0, 8'h5F, 8'h2C, 8'h37, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h35, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h30, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h45, 8'h30, 8'h37, 8'h5F, 8'h88, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'h87, 8'h5F, 8'h37, 8'h31, 8'h45, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h30, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC1, 8'h31, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h1F, 8'h39, 8'hA0, 8'hB9, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hB8, 8'hA0, 8'h39, 8'h20, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h31, 8'hC1, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hB0, 8'h31, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h43, 8'h18, 8'h40, 8'hD5, 8'hE0, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE0, 8'hD5, 8'h40, 8'h1A, 8'h43, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h31, 8'hAF, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h9B, 8'h34, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h3B, 8'h2A, 8'h5A, 8'hF6, 8'hF8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF8, 8'hF6, 8'h5A, 8'h2C, 8'h3B, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h34, 8'h9B, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD6, 8'h87, 8'h37, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h40, 8'h2C, 8'h54, 8'h83, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h83, 8'h56, 8'h2C, 8'h40, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h37, 8'h86, 8'hD6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDA, 8'h70, 8'h3B, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h3A, 8'h1A, 8'h8B, 8'hB6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB6, 8'h8B, 8'h1A, 8'h3A, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h6F, 8'hDA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDD, 8'h5D, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h36, 8'h15, 8'hB8, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hB9, 8'h15, 8'h36, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h5B, 8'hDD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDD, 8'h4C, 8'h41, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h42, 8'h35, 8'h2C, 8'hD8, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD8, 8'h2C, 8'h35, 8'h42, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h42, 8'h4B, 8'hDD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'h40, 8'h42, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3A, 8'h35, 8'h5F, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'h5F, 8'h35, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h3F, 8'hDC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h36, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h48, 8'h30, 8'h37, 8'hA0, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hA0, 8'h36, 8'h30, 8'h48, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h35, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h2E, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h2B, 8'h3F, 8'hD5, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hD5, 8'h3E, 8'h2B, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2D, 8'hD4, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCA, 8'h2B, 8'h44, 8'h45, 8'h45, 8'h45, 8'h46, 8'h41, 8'h30, 8'h59, 8'hF6, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF6, 8'h58, 8'h30, 8'h41, 8'h46, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2B, 8'hCA, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hBC, 8'h2E, 8'h44, 8'h45, 8'h45, 8'h45, 8'h46, 8'h37, 8'h3E, 8'h83, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h82, 8'h3E, 8'h37, 8'h46, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2E, 8'hBB, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hAB, 8'h33, 8'h45, 8'h45, 8'h45, 8'h45, 8'h48, 8'h2B, 8'h52, 8'hB5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hB5, 8'h52, 8'h2B, 8'h48, 8'h45, 8'h45, 8'h45, 8'h45, 8'h33, 8'hAB, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'h9C, 8'h38, 8'h45, 8'h45, 8'h45, 8'h45, 8'h47, 8'h24, 8'h67, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'h67, 8'h24, 8'h47, 8'h45, 8'h45, 8'h45, 8'h45, 8'h38, 8'h9B, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h8F, 8'h3B, 8'h45, 8'h45, 8'h45, 8'h45, 8'h42, 8'h2B, 8'h83, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'h83, 8'h2B, 8'h42, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3B, 8'h8E, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h85, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3A, 8'h3E, 8'hA4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hA4, 8'h3E, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h84, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h7B, 8'h3D, 8'h45, 8'h45, 8'h45, 8'h46, 8'h30, 8'h57, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'h57, 8'h30, 8'h46, 8'h45, 8'h45, 8'h45, 8'h3D, 8'h7B, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h72, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h46, 8'h29, 8'h70, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFB, 8'hFA, 8'hF9, 8'hF8, 8'hF7, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF6, 8'hF7, 8'hF8, 8'hF9, 8'hFA, 8'hFB, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'h70, 8'h29, 8'h46, 8'h45, 8'h45, 8'h45, 8'h3E, 8'h72, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD6, 8'h6A, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h43, 8'h2B, 8'h8E, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF4, 8'hED, 8'hE8, 8'hE3, 8'hDE, 8'hDA, 8'hD6, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD5, 8'hD6, 8'hDA, 8'hDE, 8'hE3, 8'hE8, 8'hED, 8'hF4, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'h8E, 8'h2B, 8'h43, 8'h45, 8'h45, 8'h45, 8'h3E, 8'h6A, 8'hD6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD7, 8'h62, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h35, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hE6, 8'hD7, 8'hCA, 8'hBE, 8'hB4, 8'hAA, 8'hA2, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA0, 8'hA2, 8'hAB, 8'hB5, 8'hBE, 8'hCB, 8'hD7, 8'hE6, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h35, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h62, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h5B, 8'h40, 8'h45, 8'h45, 8'h45, 8'h3A, 8'h42, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hD5, 8'hBC, 8'hA6, 8'h92, 8'h80, 8'h70, 8'h63, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h5F, 8'h62, 8'h71, 8'h81, 8'h92, 8'hA8, 8'hBC, 8'hD6, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'h42, 8'h3A, 8'h45, 8'h45, 8'h45, 8'h40, 8'h5B, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h54, 8'h41, 8'h45, 8'h45, 8'h45, 8'h36, 8'h53, 8'hEA, 8'hFE, 8'hFB, 8'hF9, 8'hF7, 8'hF6, 8'hF6, 8'hE1, 8'hC1, 8'hA1, 8'h86, 8'h6C, 8'h56, 8'h42, 8'h31, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h2C, 8'h30, 8'h43, 8'h58, 8'h6C, 8'h88, 8'hA1, 8'hC2, 8'hE2, 8'hF6, 8'hF6, 8'hF7, 8'hF9, 8'hFB, 8'hFE, 8'hEA, 8'h53, 8'h36, 8'h45, 8'h45, 8'h45, 8'h41, 8'h54, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h4E, 8'h41, 8'h45, 8'h45, 8'h44, 8'h36, 8'h70, 8'hFA, 8'hFA, 8'hEE, 8'hE4, 8'hDA, 8'hD5, 8'hD5, 8'hC2, 8'hA3, 8'h85, 8'h6A, 8'h52, 8'h3D, 8'h29, 8'h19, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h18, 8'h2B, 8'h3E, 8'h52, 8'h6D, 8'h85, 8'hA4, 8'hC3, 8'hD5, 8'hD5, 8'hDA, 8'hE4, 8'hEE, 8'hFA, 8'hFA, 8'h70, 8'h36, 8'h44, 8'h45, 8'h45, 8'h41, 8'h4E, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD0, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDA, 8'h4A, 8'h42, 8'h45, 8'h45, 8'h44, 8'h3A, 8'h95, 8'hFF, 8'hF4, 8'hD9, 8'hC1, 8'hAA, 8'hA0, 8'hA0, 8'h94, 8'h7E, 8'h69, 8'h56, 8'h45, 8'h36, 8'h28, 8'h1D, 8'h1B, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1B, 8'h1D, 8'h2A, 8'h37, 8'h45, 8'h58, 8'h69, 8'h7E, 8'h94, 8'hA0, 8'hA0, 8'hAA, 8'hC1, 8'hD9, 8'hF4, 8'hFF, 8'h95, 8'h3A, 8'h44, 8'h45, 8'h45, 8'h42, 8'h4A, 8'hDA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDA, 8'h45, 8'h42, 8'h45, 8'h45, 8'h42, 8'h40, 8'hC0, 8'hFF, 8'hED, 8'hC0, 8'h96, 8'h6F, 8'h5F, 8'h5F, 8'h5C, 8'h53, 8'h4B, 8'h43, 8'h3D, 8'h37, 8'h32, 8'h2D, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2E, 8'h2D, 8'h32, 8'h38, 8'h3D, 8'h44, 8'h4B, 8'h53, 8'h5D, 8'h5F, 8'h5F, 8'h6F, 8'h96, 8'hC0, 8'hED, 8'hFF, 8'hC0, 8'h40, 8'h42, 8'h45, 8'h45, 8'h42, 8'h45, 8'hDA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h42, 8'h43, 8'h45, 8'h45, 8'h42, 8'h47, 8'hDC, 8'hF6, 8'hDF, 8'hA6, 8'h72, 8'h41, 8'h2C, 8'h2C, 8'h31, 8'h32, 8'h34, 8'h35, 8'h37, 8'h38, 8'h39, 8'h3A, 8'h3D, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3E, 8'h3D, 8'h3B, 8'h3A, 8'h38, 8'h37, 8'h36, 8'h34, 8'h32, 8'h31, 8'h2C, 8'h2C, 8'h41, 8'h72, 8'hA6, 8'hDF, 8'hF6, 8'hDC, 8'h47, 8'h42, 8'h45, 8'h45, 8'h43, 8'h42, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3E, 8'h43, 8'h45, 8'h45, 8'h41, 8'h52, 8'hD6, 8'hD5, 8'hC0, 8'h8A, 8'h57, 8'h28, 8'h15, 8'h15, 8'h1D, 8'h23, 8'h2B, 8'h30, 8'h36, 8'h3A, 8'h3F, 8'h42, 8'h46, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h46, 8'h43, 8'h3F, 8'h3A, 8'h36, 8'h30, 8'h2B, 8'h23, 8'h1D, 8'h15, 8'h15, 8'h28, 8'h57, 8'h89, 8'hC0, 8'hD5, 8'hD6, 8'h52, 8'h41, 8'h45, 8'h45, 8'h43, 8'h3E, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3C, 8'h43, 8'h45, 8'h45, 8'h40, 8'h60, 8'hAF, 8'hA0, 8'h92, 8'h6C, 8'h49, 8'h28, 8'h1B, 8'h1C, 8'h22, 8'h28, 8'h2F, 8'h34, 8'h39, 8'h3D, 8'h41, 8'h44, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h45, 8'h41, 8'h3D, 8'h39, 8'h34, 8'h2F, 8'h27, 8'h22, 8'h1C, 8'h1B, 8'h28, 8'h49, 8'h6B, 8'h92, 8'hA0, 8'hB0, 8'h61, 8'h40, 8'h45, 8'h45, 8'h43, 8'h3C, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3B, 8'h44, 8'h45, 8'h45, 8'h3F, 8'h71, 8'h79, 8'h5F, 8'h5B, 8'h4D, 8'h3E, 8'h32, 8'h2E, 8'h2E, 8'h32, 8'h35, 8'h38, 8'h3B, 8'h3E, 8'h41, 8'h43, 8'h45, 8'h46, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h46, 8'h45, 8'h43, 8'h41, 8'h3E, 8'h3B, 8'h38, 8'h35, 8'h32, 8'h2E, 8'h2E, 8'h32, 8'h3E, 8'h4C, 8'h5B, 8'h5F, 8'h7A, 8'h71, 8'h3F, 8'h45, 8'h45, 8'h44, 8'h3B, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h39, 8'h44, 8'h45, 8'h45, 8'h3F, 8'h7B, 8'h4D, 8'h2C, 8'h30, 8'h35, 8'h37, 8'h3A, 8'h3D, 8'h3E, 8'h3F, 8'h40, 8'h41, 8'h42, 8'h43, 8'h44, 8'h44, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h44, 8'h44, 8'h43, 8'h42, 8'h41, 8'h3F, 8'h3F, 8'h3E, 8'h3D, 8'h3A, 8'h37, 8'h33, 8'h30, 8'h2C, 8'h4E, 8'h7C, 8'h3F, 8'h45, 8'h45, 8'h44, 8'h39, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h39, 8'h44, 8'h45, 8'h45, 8'h3F, 8'h78, 8'h34, 8'h15, 8'h1D, 8'h2A, 8'h34, 8'h3F, 8'h46, 8'h47, 8'h46, 8'h46, 8'h45, 8'h46, 8'h45, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h46, 8'h45, 8'h46, 8'h45, 8'h46, 8'h46, 8'h47, 8'h46, 8'h3F, 8'h34, 8'h29, 8'h1D, 8'h15, 8'h35, 8'h79, 8'h3F, 8'h45, 8'h45, 8'h44, 8'h39, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3B, 8'h44, 8'h45, 8'h45, 8'h41, 8'h69, 8'h30, 8'h1B, 8'h22, 8'h2E, 8'h38, 8'h42, 8'h48, 8'h48, 8'h48, 8'h47, 8'h46, 8'h47, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h47, 8'h46, 8'h47, 8'h48, 8'h48, 8'h48, 8'h42, 8'h38, 8'h2D, 8'h22, 8'h1B, 8'h31, 8'h69, 8'h41, 8'h45, 8'h45, 8'h44, 8'h3B, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3C, 8'h43, 8'h45, 8'h45, 8'h43, 8'h52, 8'h35, 8'h2E, 8'h32, 8'h38, 8'h3D, 8'h43, 8'h46, 8'h47, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h47, 8'h46, 8'h46, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h48, 8'h48, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h47, 8'h46, 8'h46, 8'h47, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h47, 8'h46, 8'h43, 8'h3D, 8'h38, 8'h32, 8'h2E, 8'h35, 8'h52, 8'h43, 8'h45, 8'h45, 8'h43, 8'h3C, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3F, 8'h43, 8'h45, 8'h45, 8'h45, 8'h41, 8'h39, 8'h3D, 8'h3F, 8'h40, 8'h42, 8'h44, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h46, 8'h45, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h46, 8'h45, 8'h46, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h44, 8'h42, 8'h41, 8'h3F, 8'h3D, 8'h39, 8'h40, 8'h45, 8'h45, 8'h45, 8'h43, 8'h3F, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h43, 8'h43, 8'h45, 8'h45, 8'h46, 8'h38, 8'h3D, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h45, 8'h44, 8'h43, 8'h42, 8'h42, 8'h41, 8'h40, 8'h40, 8'h40, 8'h3F, 8'h3F, 8'h3E, 8'h3E, 8'h3F, 8'h3F, 8'h3E, 8'h3E, 8'h3F, 8'h3F, 8'h40, 8'h40, 8'h40, 8'h41, 8'h42, 8'h42, 8'h43, 8'h44, 8'h45, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h3C, 8'h38, 8'h46, 8'h45, 8'h45, 8'h43, 8'h43, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDA, 8'h48, 8'h42, 8'h45, 8'h45, 8'h46, 8'h39, 8'h40, 8'h48, 8'h48, 8'h46, 8'h46, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h42, 8'h40, 8'h3D, 8'h3C, 8'h39, 8'h38, 8'h37, 8'h35, 8'h34, 8'h33, 8'h32, 8'h32, 8'h32, 8'h32, 8'h32, 8'h32, 8'h33, 8'h34, 8'h35, 8'h37, 8'h38, 8'h39, 8'h3C, 8'h3D, 8'h40, 8'h42, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h46, 8'h47, 8'h48, 8'h48, 8'h3F, 8'h39, 8'h46, 8'h45, 8'h45, 8'h42, 8'h48, 8'hDA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE1, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h4E, 8'h42, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h42, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h47, 8'h48, 8'h46, 8'h41, 8'h3C, 8'h38, 8'h34, 8'h30, 8'h2D, 8'h2A, 8'h28, 8'h26, 8'h24, 8'h24, 8'h23, 8'h22, 8'h22, 8'h23, 8'h24, 8'h24, 8'h26, 8'h28, 8'h2A, 8'h2D, 8'h30, 8'h34, 8'h38, 8'h3C, 8'h41, 8'h46, 8'h48, 8'h47, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h42, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h42, 8'h4E, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h55, 8'h41, 8'h45, 8'h45, 8'h45, 8'h43, 8'h44, 8'h46, 8'h46, 8'h45, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h44, 8'h3E, 8'h39, 8'h35, 8'h31, 8'h2C, 8'h2A, 8'h27, 8'h24, 8'h22, 8'h20, 8'h1F, 8'h1F, 8'h1D, 8'h1D, 8'h1F, 8'h1F, 8'h20, 8'h22, 8'h24, 8'h27, 8'h2A, 8'h2C, 8'h31, 8'h35, 8'h39, 8'h3E, 8'h44, 8'h46, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h44, 8'h43, 8'h45, 8'h45, 8'h45, 8'h41, 8'h55, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD7, 8'h61, 8'h3D, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h45, 8'h44, 8'h42, 8'h41, 8'h40, 8'h3F, 8'h3D, 8'h3B, 8'h3A, 8'h39, 8'h38, 8'h37, 8'h37, 8'h35, 8'h35, 8'h34, 8'h33, 8'h34, 8'h34, 8'h32, 8'h32, 8'h34, 8'h34, 8'h33, 8'h34, 8'h35, 8'h35, 8'h37, 8'h36, 8'h38, 8'h39, 8'h3A, 8'h3B, 8'h3D, 8'h3F, 8'h40, 8'h41, 8'h42, 8'h44, 8'h45, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3D, 8'h61, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD6, 8'h6F, 8'h39, 8'h46, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h41, 8'h3D, 8'h39, 8'h36, 8'h32, 8'h30, 8'h37, 8'h3D, 8'h44, 8'h49, 8'h4E, 8'h52, 8'h56, 8'h59, 8'h5B, 8'h5D, 8'h5F, 8'h60, 8'h5F, 8'h5F, 8'h60, 8'h5F, 8'h5D, 8'h5B, 8'h59, 8'h56, 8'h52, 8'h4E, 8'h49, 8'h43, 8'h3D, 8'h37, 8'h30, 8'h32, 8'h36, 8'h39, 8'h3D, 8'h41, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h46, 8'h39, 8'h6F, 8'hD6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h80, 8'h33, 8'h47, 8'h46, 8'h46, 8'h46, 8'h47, 8'h47, 8'h48, 8'h46, 8'h3E, 8'h36, 8'h30, 8'h29, 8'h23, 8'h21, 8'h32, 8'h43, 8'h52, 8'h60, 8'h6D, 8'h77, 8'h7F, 8'h88, 8'h8E, 8'h92, 8'h97, 8'h99, 8'h99, 8'h99, 8'h99, 8'h97, 8'h92, 8'h8E, 8'h88, 8'h7F, 8'h77, 8'h6B, 8'h60, 8'h52, 8'h43, 8'h32, 8'h20, 8'h23, 8'h29, 8'h30, 8'h36, 8'h3E, 8'h46, 8'h48, 8'h47, 8'h47, 8'h46, 8'h46, 8'h46, 8'h47, 8'h33, 8'h7F, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h90, 8'h2F, 8'h46, 8'h45, 8'h45, 8'h45, 8'h46, 8'h46, 8'h46, 8'h44, 8'h3B, 8'h33, 8'h2C, 8'h25, 8'h1E, 8'h1D, 8'h36, 8'h4D, 8'h63, 8'h76, 8'h88, 8'h96, 8'hA2, 8'hAE, 8'hB7, 8'hBD, 8'hC3, 8'hC6, 8'hC8, 8'hC8, 8'hC6, 8'hC3, 8'hBD, 8'hB7, 8'hAE, 8'hA2, 8'h96, 8'h87, 8'h76, 8'h62, 8'h4D, 8'h36, 8'h1C, 8'h1E, 8'h25, 8'h2C, 8'h33, 8'h3B, 8'h44, 8'h46, 8'h46, 8'h46, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2F, 8'h90, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'hA4, 8'h2F, 8'h41, 8'h44, 8'h44, 8'h43, 8'h42, 8'h40, 8'h3F, 8'h3D, 8'h3B, 8'h39, 8'h37, 8'h35, 8'h33, 8'h34, 8'h4E, 8'h66, 8'h7C, 8'h8E, 8'hA1, 8'hAF, 8'hBB, 8'hC7, 8'hCF, 8'hD6, 8'hDC, 8'hDF, 8'hE1, 8'hE1, 8'hDF, 8'hDC, 8'hD6, 8'hCF, 8'hC7, 8'hBB, 8'hAF, 8'hA0, 8'h8E, 8'h7B, 8'h66, 8'h4E, 8'h34, 8'h33, 8'h35, 8'h37, 8'h39, 8'h3B, 8'h3D, 8'h3F, 8'h40, 8'h42, 8'h43, 8'h44, 8'h44, 8'h41, 8'h2F, 8'hA3, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hB8, 8'h32, 8'h38, 8'h41, 8'h42, 8'h3F, 8'h3B, 8'h37, 8'h32, 8'h32, 8'h3C, 8'h46, 8'h4F, 8'h57, 8'h5F, 8'h65, 8'h7A, 8'h8B, 8'h9A, 8'hA7, 8'hB5, 8'hBF, 8'hC8, 8'hD0, 8'hD6, 8'hDA, 8'hDF, 8'hE1, 8'hE2, 8'hE2, 8'hE1, 8'hDF, 8'hDA, 8'hD6, 8'hD0, 8'hC8, 8'hBF, 8'hB4, 8'hA7, 8'h9A, 8'h8B, 8'h7A, 8'h65, 8'h5F, 8'h57, 8'h4F, 8'h46, 8'h3C, 8'h31, 8'h32, 8'h37, 8'h3B, 8'h3F, 8'h42, 8'h41, 8'h38, 8'h32, 8'hB8, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCF, 8'h37, 8'h2E, 8'h3D, 8'h40, 8'h3B, 8'h33, 8'h2B, 8'h23, 8'h24, 8'h3F, 8'h56, 8'h6D, 8'h83, 8'h98, 8'hA4, 8'hB0, 8'hB8, 8'hBE, 8'hC3, 8'hC8, 8'hCC, 8'hD0, 8'hD4, 8'hD5, 8'hD7, 8'hD9, 8'hD9, 8'hDA, 8'hDA, 8'hD9, 8'hD9, 8'hD7, 8'hD5, 8'hD4, 8'hD0, 8'hCC, 8'hC8, 8'hC3, 8'hBD, 8'hB8, 8'hB0, 8'hA3, 8'h98, 8'h83, 8'h6D, 8'h56, 8'h3D, 8'h23, 8'h23, 8'h2B, 8'h33, 8'h3B, 8'h40, 8'h3D, 8'h2E, 8'h37, 8'hCE, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDF, 8'h42, 8'h29, 8'h3B, 8'h3D, 8'h38, 8'h30, 8'h27, 8'h1E, 8'h21, 8'h47, 8'h69, 8'h89, 8'hA8, 8'hC5, 8'hD5, 8'hDA, 8'hDB, 8'hD9, 8'hD7, 8'hD7, 8'hD7, 8'hD6, 8'hD6, 8'hD4, 8'hD3, 8'hD4, 8'hD3, 8'hD3, 8'hD3, 8'hD3, 8'hD4, 8'hD3, 8'hD4, 8'hD6, 8'hD6, 8'hD7, 8'hD7, 8'hD7, 8'hD9, 8'hDB, 8'hDA, 8'hD5, 8'hC5, 8'hA8, 8'h89, 8'h69, 8'h46, 8'h20, 8'h1E, 8'h27, 8'h30, 8'h38, 8'h3D, 8'h3B, 8'h29, 8'h42, 8'hDF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE5, 8'h5D, 8'h32, 8'h3A, 8'h3A, 8'h3A, 8'h38, 8'h36, 8'h32, 8'h39, 8'h60, 8'h82, 8'hA2, 8'hC0, 8'hDF, 8'hED, 8'hEE, 8'hEB, 8'hE5, 8'hE1, 8'hDD, 8'hDA, 8'hD8, 8'hD5, 8'hD3, 8'hD1, 8'hD0, 8'hCF, 8'hCF, 8'hCF, 8'hCF, 8'hD0, 8'hD1, 8'hD3, 8'hD5, 8'hD8, 8'hDA, 8'hDE, 8'hE1, 8'hE5, 8'hEB, 8'hEE, 8'hED, 8'hDF, 8'hC0, 8'hA2, 8'h82, 8'h5F, 8'h37, 8'h32, 8'h35, 8'h38, 8'h3A, 8'h3A, 8'h3A, 8'h32, 8'h5D, 8'hE5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE0, 8'h85, 8'h49, 8'h3B, 8'h38, 8'h3F, 8'h4A, 8'h55, 8'h5E, 8'h69, 8'h87, 8'h9F, 8'hB6, 8'hCB, 8'hE1, 8'hEB, 8'hEB, 8'hE7, 8'hE2, 8'hDE, 8'hDA, 8'hD8, 8'hD5, 8'hD3, 8'hD1, 8'hCF, 8'hCE, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCE, 8'hCF, 8'hD1, 8'hD3, 8'hD5, 8'hD8, 8'hDB, 8'hDE, 8'hE2, 8'hE7, 8'hEB, 8'hEB, 8'hE1, 8'hCB, 8'hB6, 8'h9F, 8'h86, 8'h68, 8'h5E, 8'h54, 8'h4A, 8'h3F, 8'h38, 8'h3B, 8'h49, 8'h85, 8'hE0, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD7, 8'hB7, 8'h66, 8'h3C, 8'h34, 8'h47, 8'h62, 8'h7D, 8'h97, 8'hA6, 8'hB6, 8'hC0, 8'hC8, 8'hD1, 8'hDA, 8'hDC, 8'hDC, 8'hDB, 8'hD8, 8'hD6, 8'hD4, 8'hD2, 8'hD1, 8'hD0, 8'hCE, 8'hCD, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCD, 8'hCE, 8'hD0, 8'hD1, 8'hD2, 8'hD4, 8'hD6, 8'hD8, 8'hDB, 8'hDC, 8'hDC, 8'hDA, 8'hD1, 8'hC8, 8'hC0, 8'hB6, 8'hA5, 8'h97, 8'h7C, 8'h62, 8'h47, 8'h34, 8'h3C, 8'h66, 8'hB7, 8'hD7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hDD, 8'h81, 8'h45, 8'h39, 8'h53, 8'h79, 8'h9F, 8'hC4, 8'hD6, 8'hDB, 8'hD9, 8'hD7, 8'hD5, 8'hD4, 8'hD1, 8'hD1, 8'hD1, 8'hD0, 8'hCF, 8'hCE, 8'hCE, 8'hCD, 8'hCD, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCD, 8'hCD, 8'hCE, 8'hCE, 8'hCF, 8'hD0, 8'hD1, 8'hD1, 8'hD1, 8'hD4, 8'hD5, 8'hD7, 8'hD9, 8'hDB, 8'hD6, 8'hC4, 8'h9E, 8'h79, 8'h53, 8'h39, 8'h45, 8'h81, 8'hDD, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hEE, 8'h9B, 8'h5D, 8'h52, 8'h6C, 8'h92, 8'hB8, 8'hDD, 8'hED, 8'hEC, 8'hE5, 8'hDD, 8'hD6, 8'hD0, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hD0, 8'hD6, 8'hDD, 8'hE5, 8'hED, 8'hED, 8'hDD, 8'hB7, 8'h92, 8'h6C, 8'h52, 8'h5D, 8'h9B, 8'hEE, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hEA, 8'hB1, 8'h85, 8'h7D, 8'h8F, 8'hAA, 8'hC5, 8'hE0, 8'hEA, 8'hE8, 8'hE1, 8'hDA, 8'hD4, 8'hCE, 8'hC9, 8'hC9, 8'hCA, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCA, 8'hCA, 8'hC9, 8'hC9, 8'hCE, 8'hD4, 8'hDA, 8'hE1, 8'hE9, 8'hEA, 8'hE0, 8'hC5, 8'hAA, 8'h8F, 8'h7D, 8'h85, 8'hB1, 8'hEA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'hC6, 8'hB4, 8'hB1, 8'hB9, 8'hC4, 8'hCF, 8'hD9, 8'hDC, 8'hDB, 8'hD8, 8'hD4, 8'hD0, 8'hCD, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCD, 8'hD0, 8'hD4, 8'hD8, 8'hDB, 8'hDC, 8'hD9, 8'hCE, 8'hC4, 8'hB9, 8'hB1, 8'hB4, 8'hC6, 8'hDC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD1, 8'hD7, 8'hDA, 8'hDA, 8'hDA, 8'hD8, 8'hD5, 8'hD4, 8'hD0, 8'hD0, 8'hCF, 8'hCE, 8'hCD, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCD, 8'hCE, 8'hCF, 8'hD1, 8'hD0, 8'hD4, 8'hD6, 8'hD8, 8'hDA, 8'hDA, 8'hDA, 8'hD7, 8'hD1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDE, 8'hEB, 8'hEE, 8'hE9, 8'hE0, 8'hD8, 8'hD0, 8'hCA, 8'hCA, 8'hCB, 8'hCB, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCA, 8'hD0, 8'hD8, 8'hE0, 8'hE9, 8'hEE, 8'hEB, 8'hDE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDC, 8'hE8, 8'hEA, 8'hE5, 8'hDD, 8'hD5, 8'hCE, 8'hC9, 8'hC9, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCA, 8'hC9, 8'hC9, 8'hCE, 8'hD6, 8'hDD, 8'hE5, 8'hEA, 8'hE8, 8'hDC, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD4, 8'hDB, 8'hDC, 8'hDA, 8'hD6, 8'hD1, 8'hCD, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCA, 8'hCD, 8'hD1, 8'hD6, 8'hDA, 8'hDC, 8'hDB, 8'hD4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hD1, 8'hD1, 8'hD0, 8'hCF, 8'hCD, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCD, 8'hCF, 8'hD0, 8'hD1, 8'hD1, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hC9, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCA, 8'hC9, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hCD, 8'hCE, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hCE, 8'hCD, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hD1, 8'hD2, 8'hD0, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD0, 8'hD2, 8'hD1, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hCE, 8'hD6, 8'hD7, 8'hD3, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hD3, 8'hD7, 8'hD6, 8'hCE, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD0, 8'hD8, 8'hDA, 8'hD5, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD5, 8'hDA, 8'hD8, 8'hD0, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD1, 8'hD4, 8'hD5, 8'hD6, 8'hD5, 8'hD1, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hD1, 8'hD5, 8'hD6, 8'hD5, 8'hD4, 8'hD1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'hD9, 8'hCD, 8'hCB, 8'hD2, 8'hDC, 8'hD1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD1, 8'hDC, 8'hD2, 8'hCB, 8'hCD, 8'hD9, 8'hDC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF0, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hE9, 8'hE0, 8'hC2, 8'hBE, 8'hCF, 8'hEB, 8'hD7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD7, 8'hEB, 8'hCF, 8'hBE, 8'hC2, 8'hE0, 8'hE9, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hEE, 8'hDD, 8'hB4, 8'hAE, 8'hC5, 8'hED, 8'hD9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD9, 8'hED, 8'hC5, 8'hAE, 8'hB4, 8'hDD, 8'hEE, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD3, 8'hDC, 8'hC3, 8'h9B, 8'h95, 8'hAC, 8'hD6, 8'hD7, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hD7, 8'hD6, 8'hAC, 8'h95, 8'h9B, 8'hC3, 8'hDD, 8'hD3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDB, 8'hB7, 8'h95, 8'h7A, 8'h76, 8'h85, 8'hA6, 8'hCF, 8'hD3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD3, 8'hCF, 8'hA6, 8'h85, 8'h76, 8'h7A, 8'h95, 8'hB8, 8'hDB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hE5, 8'h88, 8'h5C, 8'h53, 8'h52, 8'h57, 8'h6A, 8'hC6, 8'hDB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDB, 8'hC6, 8'h6A, 8'h57, 8'h52, 8'h53, 8'h5C, 8'h89, 8'hE5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hE6, 8'h60, 8'h2F, 8'h35, 8'h36, 8'h33, 8'h3A, 8'hB7, 8'hDF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDF, 8'hB7, 8'h3A, 8'h33, 8'h36, 8'h35, 8'h2F, 8'h62, 8'hE6, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'hD0, 8'h47, 8'h1B, 8'h28, 8'h2A, 8'h22, 8'h22, 8'h9C, 8'hDC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'h9C, 8'h22, 8'h22, 8'h2A, 8'h28, 8'h1B, 8'h48, 8'hD0, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD9, 8'hA6, 8'h3D, 8'h20, 8'h2C, 8'h2D, 8'h27, 8'h24, 8'h77, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h77, 8'h24, 8'h27, 8'h2D, 8'h2C, 8'h20, 8'h3E, 8'hA5, 8'hD9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'h70, 8'h3A, 8'h30, 8'h37, 8'h38, 8'h34, 8'h31, 8'h4C, 8'hC7, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC7, 8'h4C, 8'h31, 8'h34, 8'h38, 8'h37, 8'h30, 8'h39, 8'h6F, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE5, 8'h45, 8'h38, 8'h3D, 8'h41, 8'h40, 8'h3F, 8'h3C, 8'h2A, 8'hB8, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hB8, 8'h2A, 8'h3C, 8'h3F, 8'h40, 8'h41, 8'h3D, 8'h37, 8'h44, 8'hE5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h2D, 8'h38, 8'h45, 8'h46, 8'h45, 8'h46, 8'h42, 8'h1C, 8'hA0, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'hA0, 8'h1C, 8'h42, 8'h46, 8'h45, 8'h46, 8'h45, 8'h37, 8'h2B, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC5, 8'h29, 8'h3B, 8'h47, 8'h47, 8'h46, 8'h47, 8'h44, 8'h22, 8'h80, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h80, 8'h22, 8'h44, 8'h47, 8'h46, 8'h47, 8'h47, 8'h3A, 8'h28, 8'hC5, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hAA, 8'h2E, 8'h40, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h31, 8'h5B, 8'hDF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDF, 8'h5B, 8'h31, 8'h45, 8'h46, 8'h46, 8'h46, 8'h46, 8'h40, 8'h2E, 8'hAA, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h91, 8'h32, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3D, 8'h3D, 8'hE2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE2, 8'h3D, 8'h3D, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h33, 8'h91, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h7B, 8'h37, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h2C, 8'hDD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDD, 8'h2C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h37, 8'h7B, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD7, 8'h6A, 8'h3A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2A, 8'hD2, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hD1, 8'h2A, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3B, 8'h6A, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h59, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2D, 8'hC2, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC2, 8'h2D, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3E, 8'h59, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h4B, 8'h41, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h30, 8'hB5, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hB4, 8'h30, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h41, 8'h4C, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h41, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h33, 8'hA8, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hA8, 8'h33, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h41, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h39, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h36, 8'h9E, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'h9E, 8'h36, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h3A, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCF, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h34, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h38, 8'h95, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h96, 8'h38, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h34, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h2F, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3A, 8'h8D, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8F, 8'h3A, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h30, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD7, 8'h2D, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h89, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2E, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h2E, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h88, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8A, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2F, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h31, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8A, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8A, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h31, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDC, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h33, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8A, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h33, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h34, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8B, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h34, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE1, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h34, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8B, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h34, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8C, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8C, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD0, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h34, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8B, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h34, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h34, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8B, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h34, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h33, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8B, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8B, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h33, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDE, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h31, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3C, 8'h8A, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h8A, 8'h3C, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h31, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h2E, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3B, 8'h89, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h89, 8'h3B, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2E, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD6, 8'h2D, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3B, 8'h8A, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8A, 8'h3B, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2D, 8'hD6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD8, 8'h2F, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3A, 8'h8D, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8E, 8'h3A, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h2F, 8'hD8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h33, 8'h44, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h39, 8'h94, 8'hD2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD2, 8'h94, 8'h39, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h44, 8'h33, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDA, 8'h38, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h37, 8'h9B, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'h9D, 8'h37, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h38, 8'hDA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h3F, 8'h43, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h35, 8'hA4, 8'hD0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD0, 8'hA6, 8'h35, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h43, 8'h3F, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'h49, 8'h41, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h32, 8'hB0, 8'hCF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCF, 8'hB2, 8'h32, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h41, 8'h49, 8'hDB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h56, 8'h3F, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h2E, 8'hBF, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC0, 8'h2E, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3F, 8'h56, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD7, 8'h66, 8'h3B, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h29, 8'hCF, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hD0, 8'h29, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h3B, 8'h66, 8'hD7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD5, 8'h76, 8'h38, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h2A, 8'hDC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDC, 8'h2A, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h45, 8'h38, 8'h76, 8'hD5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD3, 8'h8C, 8'h33, 8'h44, 8'h46, 8'h45, 8'h45, 8'h45, 8'h45, 8'h3E, 8'h39, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'h39, 8'h3E, 8'h45, 8'h45, 8'h45, 8'h45, 8'h46, 8'h44, 8'h33, 8'h8C, 8'hD3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'hA6, 8'h2D, 8'h41, 8'h46, 8'h46, 8'h46, 8'h46, 8'h45, 8'h33, 8'h55, 8'hDF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDF, 8'h55, 8'h33, 8'h46, 8'h46, 8'h46, 8'h46, 8'h46, 8'h41, 8'h2D, 8'hA6, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC2, 8'h25, 8'h3E, 8'h48, 8'h46, 8'h46, 8'h47, 8'h45, 8'h24, 8'h79, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h79, 8'h24, 8'h46, 8'h47, 8'h46, 8'h46, 8'h48, 8'h3E, 8'h25, 8'hC2, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD9, 8'h27, 8'h3B, 8'h46, 8'h45, 8'h45, 8'h46, 8'h43, 8'h1E, 8'h98, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'h98, 8'h1E, 8'h44, 8'h46, 8'h45, 8'h45, 8'h46, 8'h3B, 8'h27, 8'hD9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE3, 8'h3F, 8'h38, 8'h3F, 8'h40, 8'h41, 8'h40, 8'h3B, 8'h2B, 8'hB1, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'hB1, 8'h2B, 8'h3D, 8'h40, 8'h41, 8'h40, 8'h3F, 8'h38, 8'h3E, 8'hE3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'h6A, 8'h36, 8'h32, 8'h38, 8'h39, 8'h36, 8'h2F, 8'h48, 8'hC2, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hC2, 8'h48, 8'h30, 8'h36, 8'h39, 8'h38, 8'h32, 8'h36, 8'h69, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD9, 8'hA0, 8'h35, 8'h23, 8'h2E, 8'h30, 8'h2A, 8'h20, 8'h6F, 8'hD2, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hD2, 8'h6F, 8'h21, 8'h2A, 8'h30, 8'h2E, 8'h23, 8'h35, 8'h9F, 8'hD9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD3, 8'hCB, 8'h3B, 8'h1D, 8'h2A, 8'h2C, 8'h26, 8'h1C, 8'h90, 8'hDD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDD, 8'h90, 8'h1D, 8'h26, 8'h2C, 8'h2A, 8'h1D, 8'h3B, 8'hCA, 8'hD3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hE2, 8'h54, 8'h30, 8'h36, 8'h37, 8'h34, 8'h34, 8'hAB, 8'hE1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hE1, 8'hAB, 8'h34, 8'h34, 8'h37, 8'h36, 8'h30, 8'h54, 8'hE1, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hE3, 8'h7E, 8'h58, 8'h51, 8'h4F, 8'h55, 8'h65, 8'hBD, 8'hDC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'hBD, 8'h65, 8'h55, 8'h4F, 8'h51, 8'h58, 8'h7E, 8'hE2, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDB, 8'hB3, 8'h8D, 8'h72, 8'h6F, 8'h7E, 8'hA4, 8'hCC, 8'hD5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD5, 8'hCC, 8'hA4, 8'h7E, 8'h6F, 8'h72, 8'h8D, 8'hB3, 8'hDA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD8, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD4, 8'hDB, 8'hB7, 8'h90, 8'h8B, 8'hA1, 8'hD5, 8'hD7, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hD7, 8'hD5, 8'hA1, 8'h8B, 8'h90, 8'hB7, 8'hDB, 8'hD4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCF, 8'hEF, 8'hD1, 8'hA9, 8'hA3, 8'hBA, 8'hED, 8'hDC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hDC, 8'hED, 8'hBA, 8'hA3, 8'hA9, 8'hD1, 8'hEF, 8'hCF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE8, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCE, 8'hEB, 8'hD7, 8'hBB, 8'hB6, 8'hC7, 8'hEB, 8'hD9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hD9, 8'hEB, 8'hC7, 8'hB6, 8'hBB, 8'hD7, 8'hEB, 8'hCE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hE8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hDC, 8'hD6, 8'hCA, 8'hC8, 8'hCE, 8'hDD, 8'hD3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD3, 8'hDD, 8'hCE, 8'hC8, 8'hCA, 8'hD6, 8'hDC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hD1, 8'hD4, 8'hD6, 8'hD6, 8'hD4, 8'hD2, 8'hCE, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCE, 8'hD2, 8'hD4, 8'hD6, 8'hD6, 8'hD4, 8'hD1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD3, 8'hDB, 8'hDC, 8'hD6, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD6, 8'hDC, 8'hDB, 8'hD3, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hD1, 8'hD8, 8'hD9, 8'hD4, 8'hCA, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hD4, 8'hD9, 8'hD8, 8'hD1, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCE, 8'hD3, 8'hD3, 8'hD1, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hD1, 8'hD3, 8'hD3, 8'hCE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCD, 8'hCE, 8'hCE, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCE, 8'hCE, 8'hCD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hD0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hE2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC6, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCC, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hCB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD9, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hD9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEF, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hCA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC2, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC2, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC2, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hCA, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hCA, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hC1, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC1, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC2, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC2, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hC8, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC8, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE3, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hE3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEB, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC5, 8'hEB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hC6, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC6, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hCE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hCE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hC0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC0, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC6, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC6, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD4, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hD4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hBD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBD, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hC2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC2, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hCE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDD, 8'hC0, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC0, 8'hDD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hBE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBE, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hC2, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hCC, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hCC, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hD9, 8'hC1, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC1, 8'hD9, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE4, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hE4, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hC3, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC3, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hCC, 8'hC6, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC6, 8'hCC, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD7, 8'hC1, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC1, 8'hD7, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hE1, 8'hBF, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBF, 8'hE1, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hEA, 8'hC3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC3, 8'hEA, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hCC, 8'hC4, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC4, 8'hCC, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF6, 8'hD9, 8'hBF, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hBF, 8'hD9, 8'hF6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE4, 8'hBD, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBD, 8'hE4, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hED, 8'hC2, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC2, 8'hED, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hCE, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hCE, 8'hF2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hDD, 8'hBE, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBE, 8'hDD, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hEA, 8'hBB, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hBB, 8'hEA, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hF4, 8'hC2, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC2, 8'hF4, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hD1, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hD1, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hE3, 8'hBF, 8'hC9, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hC9, 8'hBF, 8'hE3, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hF3, 8'hBE, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hBE, 8'hF3, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hC4, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hC4, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC7, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC7, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE5, 8'hC5, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hC5, 8'hE5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hC7, 8'hC4, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC4, 8'hC7, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hCE, 8'hC6, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC6, 8'hCE, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'hCC, 8'hC3, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC3, 8'hCC, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hD3, 8'hBE, 8'hCB, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCB, 8'hBE, 8'hD3, 8'hE9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF5, 8'hDA, 8'hBB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hBB, 8'hDA, 8'hF5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE2, 8'hC2, 8'hC9, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC9, 8'hC2, 8'hE2, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEA, 8'hD1, 8'hC5, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hC5, 8'hD1, 8'hEA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF3, 8'hE3, 8'hC2, 8'hC5, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC5, 8'hC2, 8'hE3, 8'hF3, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF3, 8'hC1, 8'hC3, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC3, 8'hC1, 8'hF3, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hC8, 8'hC6, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC6, 8'hC8, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD5, 8'hCC, 8'hC3, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC3, 8'hCC, 8'hD5, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE6, 8'hD5, 8'hBE, 8'hC7, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC7, 8'hBE, 8'hD5, 8'hE6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDD, 8'hBB, 8'hC6, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC6, 8'hBB, 8'hDD, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hE5, 8'hC2, 8'hC6, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC6, 8'hC2, 8'hE5, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEC, 8'hD1, 8'hC8, 8'hC4, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC4, 8'hC8, 8'hD1, 8'hEC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE3, 8'hCC, 8'hBE, 8'hC8, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC8, 8'hBE, 8'hCC, 8'hE3, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hF3, 8'hD0, 8'hBC, 8'hC7, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC7, 8'hBC, 8'hD0, 8'hF3, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hD7, 8'hC3, 8'hC8, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC8, 8'hC3, 8'hD7, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE1, 8'hD1, 8'hC9, 8'hC4, 8'hC9, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hC9, 8'hC4, 8'hC9, 8'hD1, 8'hE1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hE4, 8'hCB, 8'hBE, 8'hC6, 8'hCC, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCC, 8'hC6, 8'hBE, 8'hCB, 8'hE4, 8'hEE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hF3, 8'hCE, 8'hBC, 8'hC5, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC5, 8'hBC, 8'hCE, 8'hF3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hD6, 8'hC3, 8'hC7, 8'hC8, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hC8, 8'hC7, 8'hC3, 8'hD6, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE0, 8'hD1, 8'hCB, 8'hC4, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hC4, 8'hCB, 8'hD1, 8'hE0, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hED, 8'hE4, 8'hD1, 8'hBE, 8'hC4, 8'hC9, 8'hCC, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCC, 8'hC9, 8'hC4, 8'hBE, 8'hD1, 8'hE4, 8'hED, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF7, 8'hF3, 8'hD7, 8'hBC, 8'hC2, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC2, 8'hBC, 8'hD7, 8'hF3, 8'hF7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFC, 8'hDE, 8'hC3, 8'hC6, 8'hC8, 8'hC8, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hC8, 8'hC8, 8'hC6, 8'hC3, 8'hDE, 8'hFC, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE7, 8'hD1, 8'hD0, 8'hC8, 8'hC3, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hC3, 8'hC8, 8'hD0, 8'hD1, 8'hE7, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF1, 8'hE4, 8'hDC, 8'hC9, 8'hBE, 8'hC4, 8'hC8, 8'hCB, 8'hCD, 8'hCD, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCD, 8'hCD, 8'hCB, 8'hC8, 8'hC4, 8'hBE, 8'hC9, 8'hDC, 8'hE4, 8'hF1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hF3, 8'hE7, 8'hCB, 8'hBB, 8'hC2, 8'hC7, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC7, 8'hC2, 8'hBB, 8'hCB, 8'hE7, 8'hF3, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFC, 8'hEF, 8'hD3, 8'hC2, 8'hC6, 8'hC8, 8'hC8, 8'hCA, 8'hCB, 8'hCB, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hCB, 8'hCB, 8'hC9, 8'hC8, 8'hC8, 8'hC6, 8'hC2, 8'hD3, 8'hEF, 8'hFC, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hDE, 8'hD1, 8'hCF, 8'hCA, 8'hC4, 8'hC5, 8'hC7, 8'hC9, 8'hCA, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCA, 8'hC9, 8'hC7, 8'hC5, 8'hC4, 8'hCA, 8'hCF, 8'hD1, 8'hDE, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF9, 8'hEB, 8'hE3, 8'hDC, 8'hCD, 8'hBF, 8'hC0, 8'hC4, 8'hC6, 8'hC9, 8'hCB, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCD, 8'hCB, 8'hC9, 8'hC6, 8'hC4, 8'hBF, 8'hBF, 8'hCD, 8'hDC, 8'hE3, 8'hEB, 8'hF9, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF6, 8'hF3, 8'hE6, 8'hD1, 8'hBE, 8'hBE, 8'hC2, 8'hC5, 8'hC8, 8'hCB, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCB, 8'hC8, 8'hC5, 8'hC2, 8'hBD, 8'hBE, 8'hD1, 8'hE6, 8'hF3, 8'hF6, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFC, 8'hEE, 8'hD8, 8'hC4, 8'hC4, 8'hC6, 8'hC7, 8'hC8, 8'hC8, 8'hC9, 8'hC9, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hCA, 8'hC9, 8'hC9, 8'hC9, 8'hC8, 8'hC7, 8'hC6, 8'hC4, 8'hC4, 8'hD8, 8'hEE, 8'hFC, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE2, 8'hD2, 8'hD2, 8'hCF, 8'hCC, 8'hC8, 8'hC5, 8'hC4, 8'hC5, 8'hC6, 8'hC6, 8'hC6, 8'hC7, 8'hC7, 8'hC6, 8'hC6, 8'hC6, 8'hC5, 8'hC4, 8'hC5, 8'hC8, 8'hCC, 8'hCF, 8'hD2, 8'hD2, 8'hE2, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hEE, 8'hE5, 8'hE5, 8'hDC, 8'hD2, 8'hC9, 8'hC1, 8'hBD, 8'hBF, 8'hC1, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC2, 8'hC1, 8'hBF, 8'hBD, 8'hC2, 8'hC9, 8'hD2, 8'hDC, 8'hE4, 8'hE5, 8'hEE, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF7, 8'hF3, 8'hF3, 8'hE6, 8'hD8, 8'hCB, 8'hC0, 8'hBB, 8'hBD, 8'hC0, 8'hC0, 8'hC0, 8'hC1, 8'hC1, 8'hC0, 8'hC0, 8'hC0, 8'hBD, 8'hBB, 8'hC1, 8'hCB, 8'hD8, 8'hE6, 8'hF3, 8'hF3, 8'hF7, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFC, 8'hFC, 8'hEE, 8'hE0, 8'hD3, 8'hC7, 8'hC1, 8'hC4, 8'hC6, 8'hC6, 8'hC5, 8'hC6, 8'hC6, 8'hC5, 8'hC6, 8'hC6, 8'hC4, 8'hC1, 8'hC8, 8'hD3, 8'hE0, 8'hEE, 8'hFC, 8'hFC, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF4, 8'hE8, 8'hDE, 8'hD4, 8'hD0, 8'hD2, 8'hD4, 8'hD2, 8'hD1, 8'hD0, 8'hD0, 8'hD1, 8'hD2, 8'hD4, 8'hD2, 8'hD0, 8'hD5, 8'hDE, 8'hE8, 8'hF4, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF8, 8'hF2, 8'hEB, 8'hE6, 8'hE3, 8'hE4, 8'hE5, 8'hE2, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hE2, 8'hE5, 8'hE4, 8'hE3, 8'hE6, 8'hEB, 8'hF2, 8'hF8, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFC, 8'hF9, 8'hF6, 8'hF4, 8'hF3, 8'hF3, 8'hF4, 8'hEF, 8'hEC, 8'hEA, 8'hEA, 8'hEC, 8'hEF, 8'hF4, 8'hF3, 8'hF3, 8'hF4, 8'hF6, 8'hF9, 8'hFC, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFE, 8'hFD, 8'hFD, 8'hFC, 8'hFC, 8'hFD, 8'hF8, 8'hF5, 8'hF3, 8'hF3, 8'hF5, 8'hF8, 8'hFD, 8'hFC, 8'hFC, 8'hFD, 8'hFD, 8'hFE, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hF9, 8'hF7, 8'hF7, 8'hF9, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFD, 8'hFB, 8'hFB, 8'hFB, 8'hFB, 8'hFD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFE, 8'hFD, 8'hFD, 8'hFD, 8'hFD, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF};

 reg	[7:0]	pattern_data_R2 [0:39999] = '{8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED, 8'hED}; 
 reg	[7:0]	pattern_data_B2 [0:39999] = '{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24}; 
 reg	[7:0]	pattern_data_G2 [0:39999] = '{8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C, 8'h1C};

 reg	[7:0]	pattern_data_R3 [0:39999] = '{8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F, 8'h3F}; 
 reg	[7:0]	pattern_data_B3 [0:39999] = '{8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC, 8'hCC}; 
 reg	[7:0]	pattern_data_G3 [0:39999] = '{8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48};


 reg	[7:0]	pattern_data_R4 [0:39999] = '{8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22}; 
 reg	[7:0]	pattern_data_B4 [0:39999] = '{8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C}; 
 reg	[7:0]	pattern_data_G4 [0:39999] = '{8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1, 8'hB1};
//=============================================================================
// Structural coding
//=============================================================================

					
// This signal indicate the lcd display area .
assign	display_area = ((x_cnt>(Hsync_Blank-1)&& //>215
						(x_cnt<(H_LINE-Hsync_Front_Porch))&& //< 1016
						(y_cnt>(Vertical_Back_Porch-1))&& 
						(y_cnt<(V_LINE - Vertical_Front_Porch))
						))  ? 1'b1 : 1'b0;


///////////////////////// x  y counter  and lcd hd generator //////////////////
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			x_cnt <= 11'd0;	
			mhd  <= 1'd0;  	
		end	
		else if (x_cnt == (H_LINE-1))
		begin
			x_cnt <= 11'd0;
			mhd  <= 1'd0;
		end	   
		else
		begin
			x_cnt <= x_cnt + 11'd1;
			mhd  <= 1'd1;
		end	
	end

always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
			y_cnt <= 10'd0;
		else if (x_cnt == (H_LINE-1))
		begin
			if (y_cnt == (V_LINE-1))
			begin
				y_cnt <= 10'd0;
			end
			else
				y_cnt <= y_cnt + 10'd1;	
		end
	end
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			res_cnt = 0;
			vres_cnt = 0;
		end
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin	
				if (res_cnt == (hres_limit-1))
					res_cnt = 0;	   
				else
					res_cnt = res_cnt + 1;
				if (x_cnt > (H_LINE-Hsync_Front_Porch-1))
				begin
					if (vres_cnt == (vres_limit-1))
						vres_cnt = 0;	   
					else
						vres_cnt = vres_cnt + 1;
				end
			end
		end
	end
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			res_cnt1 = 0;
			vres_cnt1 = 0;
		end
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin	
				if (res_cnt1 == (hres_limit1-1))
					res_cnt1 = 0;	   
				else
					res_cnt1 = res_cnt1 + 1;
				if (x_cnt > (H_LINE-Hsync_Front_Porch-1))
				begin
					if (vres_cnt1 == (vres_limit1-1))
						vres_cnt1 = 0;	   
					else
						vres_cnt1 = vres_cnt1 + 1;
				end
			end
		end
	end
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			pic_cnt = 99;
			pic_cnt1 = 9;
		end
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				if (res_cnt == (hres_limit - 1))
				begin
					if (pic_cnt == (0))
						pic_cnt = 99;
					else
						pic_cnt = pic_cnt - 1;
				end
				if (x_cnt > (H_LINE-Hsync_Front_Porch-1))
				begin
					if (vres_cnt ==(vres_limit-1))
					begin
						if (pic_cnt1 == tres_limit-1)
							pic_cnt1 = 9;
						else
							pic_cnt1 = pic_cnt1 + 10;
					end
					pic_cnt = pic_cnt1 + pic_cnt - 1;
				end
			end	
		end
	end

	
always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
		begin
			pic_cnt2 = 39999;
			pic_cnt3 = 99;
		end
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				if (res_cnt1 == (hres_limit1 - 1))
				begin
					if (pic_cnt2 == 0)
						pic_cnt2 = 39999;
					else
						pic_cnt2 = pic_cnt2 - 1;
				end
				if (x_cnt > (H_LINE-Hsync_Front_Porch-1))
				begin
					if (vres_cnt1 ==(vres_limit1-1))
					begin
						if (pic_cnt3 == tres_limit1-1)
							pic_cnt3 = 99;
						else
							pic_cnt3 = pic_cnt3 + 100;
					end
					pic_cnt2 = pic_cnt3 + pic_cnt2 - 1;
				end
			end	
		end
	end
////////////////////////////// touch panel timing //////////////////

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			mvd  <= 1'b1;
		else if (y_cnt == 10'd0)
			mvd  <= 1'b0;
		else
			mvd  <= 1'b1;
	end			

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			mden  <= 1'b0;
		else if (display_area)
			mden  <= 1'b1;
		else
			mden  <= 1'b0;
	end			

//////////////Picture generator ///////

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			pattern_data	<=	8'h00;
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				red_1 <= pattern_data_R1[pic_cnt2];
				green_1 <= pattern_data_G1[pic_cnt2];
				blue_1 <= pattern_data_B1[pic_cnt2];
			end
		end
end

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			pattern_data	<=	8'h00;
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				red_2 <= pattern_data_R2[pic_cnt2];
				green_2 <= pattern_data_G2[pic_cnt2];
				blue_2 <= pattern_data_B2[pic_cnt2];
			end
		end
end

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			pattern_data	<=	8'h00;
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				red_3 <= pattern_data_R3[pic_cnt2];
				green_3 <= pattern_data_G3[pic_cnt2];
				blue_3 <= pattern_data_B3[pic_cnt2];
			end
		end
end

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			pattern_data	<=	8'h00;
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch)))
		begin
			if((y_cnt>(Vertical_Back_Porch-1))&&(y_cnt<(V_LINE-Vertical_Front_Porch)))
			begin
				red_4 <= pattern_data_R4[pic_cnt2];
				green_4 <= pattern_data_G4[pic_cnt2];
				blue_4 <= pattern_data_B4[pic_cnt2];
			end
		end
end	

//////////////gray level  patten generator ///////

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			graycnt <= 0;
		else if((x_cnt>(Hsync_Blank-1))&&(x_cnt<(H_LINE-Hsync_Front_Porch))) 
			graycnt <= graycnt + 1;	
		else
			graycnt <= 0;		
end

//////////////chessboard pattern ///////

assign	msel1	=	(y_cnt>= 40 && y_cnt<88)   ?	2'b01:
						(y_cnt>=88	&& y_cnt<136)	?	2'b10	:
						(y_cnt>=136	&& y_cnt<184)	?	2'b01	:
						(y_cnt>=184	&& y_cnt<232)	?	2'b10	:
						(y_cnt>=232	&& y_cnt<280)	?	2'b01	:
						(y_cnt>=280	&& y_cnt<328)	?	2'b10	:
						(y_cnt>=328	&& y_cnt<376)	?	2'b01	:
						(y_cnt>=376	&& y_cnt<424)	?	2'b10	:
						(y_cnt>=424	&& y_cnt<472)	?	2'b01	:
						(y_cnt>=472	&& y_cnt<520)	?	2'b10	:
						   								   2'b00	;
assign	mselx1=  (x_cnt>=216 && x_cnt<296)  ?	2'b01:
						(x_cnt>=296	&& x_cnt<376)	?	2'b10	:
						(x_cnt>=376	&& x_cnt<456)	?	2'b01	:
						(x_cnt>=456	&& x_cnt<536)	?	2'b10	:
						(x_cnt>=536	&& x_cnt<616)	?	2'b01	:
						(x_cnt>=616	&& x_cnt<696)	?	2'b10	:
						(x_cnt>=696	&& x_cnt<776)	?	2'b01	:
						(x_cnt>=776	&& x_cnt<856)	?	2'b10	:
						(x_cnt>=856	&& x_cnt<936)	?	2'b01	:
						(x_cnt>=936	&& x_cnt<1016)	?	2'b10	:
						   								   2'b00	;

always@(posedge iCLK  or negedge iRST_n)
	begin
		if (!iRST_n)
			graycnt1 <= 0;
		else if(mselx1==0)
			graycnt1 <= 8'h7ff;
		else if(mselx1 ==2) 
			begin
				if(msel1 ==2)
					begin
						graycnt1 <= 8'h7f;
				end	
				else if (msel1 == 1)
					begin
						graycnt1 <= 0;
				end
				else
					graycnt1 <= 8'hff;
		end
		else if(mselx1 == 1)
				begin
				if(msel1 == 2)
					begin
						graycnt1 <= 0;
					
				end	
				else if (msel1 == 1)
					begin
						graycnt1 <= 8'h7f;						
				end
				else
					graycnt1 <= 8'hff;
		end
		else
			graycnt1 <= 0;		
end
////////////// displayed color pattern selection //////////////

assign mred    = (iDISPLAY_MODE == 2'b11)? red_2:  
				 (iDISPLAY_MODE == 2'b10)?  red_3:
			     (iDISPLAY_MODE == 2'b01)?  red_1:
										    red_4; 

assign mgreen  = (iDISPLAY_MODE == 2'b11)?  green_2: 
			     (iDISPLAY_MODE == 2'b10)?  green_3:
				 (iDISPLAY_MODE == 2'b01)?  green_1:
				  				            green_4;
				 
assign mblue   = (iDISPLAY_MODE == 2'b11)?  blue_2:  
			     (iDISPLAY_MODE == 2'b10)?  blue_3:
				 (iDISPLAY_MODE == 2'b01)?  blue_1:
				  				            blue_4;


always@(posedge iCLK or negedge iRST_n)
	begin
		if (!iRST_n)
			begin
				oHD	<= 1'd0;
				oVD	<= 1'd0;
				oDEN <= 1'd0;
				oLCD_R <= 8'd0;
				oLCD_G <= 8'd0;
				oLCD_B <= 8'd0;
			end
		else
			begin
				oHD	<= mhd;
				oVD	<= mvd;
				oDEN <= display_area;
				oLCD_R <= mred;
				oLCD_G <= mgreen;
				oLCD_B <= mblue;
			end		
	end
						
endmodule